library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity background_rom is
  port(
	  clk : in std_logic;
	  xadr: in unsigned(7 downto 0);
	  yadr : in unsigned(6 downto 0); -- 0-1023
	  rgb : out std_logic_vector(5 downto 0)
      );
end background_rom;

architecture synth of background_rom is
signal totaladr : std_logic_vector(14 downto 0);
begin
   process (clk) begin
	if rising_edge(clk) then
		case totaladr is
					when "000000000000000" => rgb <= "101111";
					when "000000000000001" => rgb <= "101111";
					when "000000000000010" => rgb <= "101111";
					when "000000000000011" => rgb <= "101111";
					when "000000000000100" => rgb <= "101111";
					when "000000000000101" => rgb <= "101111";
					when "000000000000110" => rgb <= "101111";
					when "000000000000111" => rgb <= "101111";
					when "000000000001000" => rgb <= "101111";
					when "000000000001001" => rgb <= "101111";
					when "000000000001010" => rgb <= "101111";
					when "000000000001011" => rgb <= "101111";
					when "000000000001100" => rgb <= "101111";
					when "000000000001101" => rgb <= "101111";
					when "000000000001110" => rgb <= "101111";
					when "000000000001111" => rgb <= "101111";
					when "000000000010000" => rgb <= "101111";
					when "000000000010001" => rgb <= "101111";
					when "000000000010010" => rgb <= "101111";
					when "000000000010011" => rgb <= "101111";
					when "000000000010100" => rgb <= "101111";
					when "000000000010101" => rgb <= "101111";
					when "000000000010110" => rgb <= "101111";
					when "000000000010111" => rgb <= "101111";
					when "000000000011000" => rgb <= "101111";
					when "000000000011001" => rgb <= "101111";
					when "000000000011010" => rgb <= "101111";
					when "000000000011011" => rgb <= "101111";
					when "000000000011100" => rgb <= "101111";
					when "000000000011101" => rgb <= "101111";
					when "000000000011110" => rgb <= "101111";
					when "000000000011111" => rgb <= "101111";
					when "000000000100000" => rgb <= "101111";
					when "000000000100001" => rgb <= "101111";
					when "000000000100010" => rgb <= "101111";
					when "000000000100011" => rgb <= "101111";
					when "000000000100100" => rgb <= "101111";
					when "000000000100101" => rgb <= "101111";
					when "000000000100110" => rgb <= "101111";
					when "000000000100111" => rgb <= "101111";
					when "000000000101000" => rgb <= "101111";
					when "000000000101001" => rgb <= "101111";
					when "000000000101010" => rgb <= "101111";
					when "000000000101011" => rgb <= "101111";
					when "000000000101100" => rgb <= "101111";
					when "000000000101101" => rgb <= "101111";
					when "000000000101110" => rgb <= "101111";
					when "000000000101111" => rgb <= "101111";
					when "000000000110000" => rgb <= "101111";
					when "000000000110001" => rgb <= "101111";
					when "000000000110010" => rgb <= "101111";
					when "000000000110011" => rgb <= "101111";
					when "000000000110100" => rgb <= "101111";
					when "000000000110101" => rgb <= "101111";
					when "000000000110110" => rgb <= "101111";
					when "000000000110111" => rgb <= "101111";
					when "000000000111000" => rgb <= "101111";
					when "000000000111001" => rgb <= "101111";
					when "000000000111010" => rgb <= "101111";
					when "000000000111011" => rgb <= "101111";
					when "000000000111100" => rgb <= "101111";
					when "000000000111101" => rgb <= "101111";
					when "000000000111110" => rgb <= "101111";
					when "000000000111111" => rgb <= "101111";
					when "000000001000000" => rgb <= "101111";
					when "000000001000001" => rgb <= "101111";
					when "000000001000010" => rgb <= "101111";
					when "000000001000011" => rgb <= "101111";
					when "000000001000100" => rgb <= "101111";
					when "000000001000101" => rgb <= "101111";
					when "000000001000110" => rgb <= "101111";
					when "000000001000111" => rgb <= "101111";
					when "000000001001000" => rgb <= "101111";
					when "000000001001001" => rgb <= "101111";
					when "000000001001010" => rgb <= "101111";
					when "000000001001011" => rgb <= "101111";
					when "000000001001100" => rgb <= "101111";
					when "000000001001101" => rgb <= "101111";
					when "000000001001110" => rgb <= "101111";
					when "000000001001111" => rgb <= "101111";
					when "000000001010000" => rgb <= "101111";
					when "000000001010001" => rgb <= "101111";
					when "000000001010010" => rgb <= "101111";
					when "000000001010011" => rgb <= "101111";
					when "000000001010100" => rgb <= "101111";
					when "000000001010101" => rgb <= "101111";
					when "000000001010110" => rgb <= "101111";
					when "000000001010111" => rgb <= "101111";
					when "000000001011000" => rgb <= "101111";
					when "000000001011001" => rgb <= "101111";
					when "000000001011010" => rgb <= "101111";
					when "000000001011011" => rgb <= "101111";
					when "000000001011100" => rgb <= "101111";
					when "000000001011101" => rgb <= "101111";
					when "000000001011110" => rgb <= "101111";
					when "000000001011111" => rgb <= "101111";
					when "000000001100000" => rgb <= "101111";
					when "000000001100001" => rgb <= "101111";
					when "000000001100010" => rgb <= "101111";
					when "000000001100011" => rgb <= "101111";
					when "000000001100100" => rgb <= "101111";
					when "000000001100101" => rgb <= "101111";
					when "000000001100110" => rgb <= "101111";
					when "000000001100111" => rgb <= "101111";
					when "000000001101000" => rgb <= "101111";
					when "000000001101001" => rgb <= "101111";
					when "000000001101010" => rgb <= "101111";
					when "000000001101011" => rgb <= "101111";
					when "000000001101100" => rgb <= "101111";
					when "000000001101101" => rgb <= "101111";
					when "000000001101110" => rgb <= "101111";
					when "000000001101111" => rgb <= "101111";
					when "000000001110000" => rgb <= "101111";
					when "000000001110001" => rgb <= "101111";
					when "000000001110010" => rgb <= "101111";
					when "000000001110011" => rgb <= "101111";
					when "000000001110100" => rgb <= "101111";
					when "000000001110101" => rgb <= "101111";
					when "000000001110110" => rgb <= "101111";
					when "000000001110111" => rgb <= "101111";
					when "000000001111000" => rgb <= "101111";
					when "000000001111001" => rgb <= "101111";
					when "000000001111010" => rgb <= "101111";
					when "000000001111011" => rgb <= "101111";
					when "000000001111100" => rgb <= "101111";
					when "000000001111101" => rgb <= "101111";
					when "000000001111110" => rgb <= "101111";
					when "000000001111111" => rgb <= "101111";
					when "000000010000000" => rgb <= "101111";
					when "000000010000001" => rgb <= "101111";
					when "000000010000010" => rgb <= "101111";
					when "000000010000011" => rgb <= "101111";
					when "000000010000100" => rgb <= "101111";
					when "000000010000101" => rgb <= "101111";
					when "000000010000110" => rgb <= "101111";
					when "000000010000111" => rgb <= "101111";
					when "000000010001000" => rgb <= "101111";
					when "000000010001001" => rgb <= "101111";
					when "000000010001010" => rgb <= "101111";
					when "000000010001011" => rgb <= "101111";
					when "000000010001100" => rgb <= "101111";
					when "000000010001101" => rgb <= "101111";
					when "000000010001110" => rgb <= "101111";
					when "000000010001111" => rgb <= "101111";
					when "000000010010000" => rgb <= "101111";
					when "000000010010001" => rgb <= "101111";
					when "000000010010010" => rgb <= "101111";
					when "000000010010011" => rgb <= "101111";
					when "000000010010100" => rgb <= "101111";
					when "000000010010101" => rgb <= "101111";
					when "000000010010110" => rgb <= "101111";
					when "000000010010111" => rgb <= "101111";
					when "000000010011000" => rgb <= "101111";
					when "000000010011001" => rgb <= "101111";
					when "000000010011010" => rgb <= "101111";
					when "000000010011011" => rgb <= "101111";
					when "000000010011100" => rgb <= "101111";
					when "000000010011101" => rgb <= "101111";
					when "000000010011110" => rgb <= "101111";
					when "000000010011111" => rgb <= "101111";
					when "000000100000000" => rgb <= "101111";
					when "000000100000001" => rgb <= "101111";
					when "000000100000010" => rgb <= "101111";
					when "000000100000011" => rgb <= "101111";
					when "000000100000100" => rgb <= "101111";
					when "000000100000101" => rgb <= "101111";
					when "000000100000110" => rgb <= "101111";
					when "000000100000111" => rgb <= "101111";
					when "000000100001000" => rgb <= "101111";
					when "000000100001001" => rgb <= "101111";
					when "000000100001010" => rgb <= "101111";
					when "000000100001011" => rgb <= "101111";
					when "000000100001100" => rgb <= "101111";
					when "000000100001101" => rgb <= "101111";
					when "000000100001110" => rgb <= "101111";
					when "000000100001111" => rgb <= "101111";
					when "000000100010000" => rgb <= "101111";
					when "000000100010001" => rgb <= "101111";
					when "000000100010010" => rgb <= "101111";
					when "000000100010011" => rgb <= "101111";
					when "000000100010100" => rgb <= "101111";
					when "000000100010101" => rgb <= "101111";
					when "000000100010110" => rgb <= "101111";
					when "000000100010111" => rgb <= "101111";
					when "000000100011000" => rgb <= "101111";
					when "000000100011001" => rgb <= "101111";
					when "000000100011010" => rgb <= "101111";
					when "000000100011011" => rgb <= "101111";
					when "000000100011100" => rgb <= "101111";
					when "000000100011101" => rgb <= "101111";
					when "000000100011110" => rgb <= "101111";
					when "000000100011111" => rgb <= "101111";
					when "000000100100000" => rgb <= "101111";
					when "000000100100001" => rgb <= "101111";
					when "000000100100010" => rgb <= "101111";
					when "000000100100011" => rgb <= "101111";
					when "000000100100100" => rgb <= "101111";
					when "000000100100101" => rgb <= "101111";
					when "000000100100110" => rgb <= "101111";
					when "000000100100111" => rgb <= "101111";
					when "000000100101000" => rgb <= "101111";
					when "000000100101001" => rgb <= "101111";
					when "000000100101010" => rgb <= "101111";
					when "000000100101011" => rgb <= "101111";
					when "000000100101100" => rgb <= "101111";
					when "000000100101101" => rgb <= "101111";
					when "000000100101110" => rgb <= "101111";
					when "000000100101111" => rgb <= "101111";
					when "000000100110000" => rgb <= "101111";
					when "000000100110001" => rgb <= "101111";
					when "000000100110010" => rgb <= "101111";
					when "000000100110011" => rgb <= "101111";
					when "000000100110100" => rgb <= "101111";
					when "000000100110101" => rgb <= "101111";
					when "000000100110110" => rgb <= "101111";
					when "000000100110111" => rgb <= "101111";
					when "000000100111000" => rgb <= "101111";
					when "000000100111001" => rgb <= "101111";
					when "000000100111010" => rgb <= "101111";
					when "000000100111011" => rgb <= "101111";
					when "000000100111100" => rgb <= "101111";
					when "000000100111101" => rgb <= "101111";
					when "000000100111110" => rgb <= "101111";
					when "000000100111111" => rgb <= "101111";
					when "000000101000000" => rgb <= "101111";
					when "000000101000001" => rgb <= "101111";
					when "000000101000010" => rgb <= "101111";
					when "000000101000011" => rgb <= "101111";
					when "000000101000100" => rgb <= "101111";
					when "000000101000101" => rgb <= "101111";
					when "000000101000110" => rgb <= "101111";
					when "000000101000111" => rgb <= "101111";
					when "000000101001000" => rgb <= "101111";
					when "000000101001001" => rgb <= "101111";
					when "000000101001010" => rgb <= "101111";
					when "000000101001011" => rgb <= "101111";
					when "000000101001100" => rgb <= "101111";
					when "000000101001101" => rgb <= "101111";
					when "000000101001110" => rgb <= "101111";
					when "000000101001111" => rgb <= "101111";
					when "000000101010000" => rgb <= "101111";
					when "000000101010001" => rgb <= "101111";
					when "000000101010010" => rgb <= "101111";
					when "000000101010011" => rgb <= "101111";
					when "000000101010100" => rgb <= "101111";
					when "000000101010101" => rgb <= "101111";
					when "000000101010110" => rgb <= "101111";
					when "000000101010111" => rgb <= "101111";
					when "000000101011000" => rgb <= "101111";
					when "000000101011001" => rgb <= "101111";
					when "000000101011010" => rgb <= "101111";
					when "000000101011011" => rgb <= "101111";
					when "000000101011100" => rgb <= "101111";
					when "000000101011101" => rgb <= "101111";
					when "000000101011110" => rgb <= "101111";
					when "000000101011111" => rgb <= "101111";
					when "000000101100000" => rgb <= "101111";
					when "000000101100001" => rgb <= "101111";
					when "000000101100010" => rgb <= "101111";
					when "000000101100011" => rgb <= "101111";
					when "000000101100100" => rgb <= "101111";
					when "000000101100101" => rgb <= "101111";
					when "000000101100110" => rgb <= "101111";
					when "000000101100111" => rgb <= "101111";
					when "000000101101000" => rgb <= "101111";
					when "000000101101001" => rgb <= "101111";
					when "000000101101010" => rgb <= "101111";
					when "000000101101011" => rgb <= "101111";
					when "000000101101100" => rgb <= "101111";
					when "000000101101101" => rgb <= "101111";
					when "000000101101110" => rgb <= "101111";
					when "000000101101111" => rgb <= "101111";
					when "000000101110000" => rgb <= "101111";
					when "000000101110001" => rgb <= "101111";
					when "000000101110010" => rgb <= "101111";
					when "000000101110011" => rgb <= "101111";
					when "000000101110100" => rgb <= "101111";
					when "000000101110101" => rgb <= "101111";
					when "000000101110110" => rgb <= "101111";
					when "000000101110111" => rgb <= "101111";
					when "000000101111000" => rgb <= "101111";
					when "000000101111001" => rgb <= "101111";
					when "000000101111010" => rgb <= "101111";
					when "000000101111011" => rgb <= "101111";
					when "000000101111100" => rgb <= "101111";
					when "000000101111101" => rgb <= "101111";
					when "000000101111110" => rgb <= "101111";
					when "000000101111111" => rgb <= "101111";
					when "000000110000000" => rgb <= "101111";
					when "000000110000001" => rgb <= "101111";
					when "000000110000010" => rgb <= "101111";
					when "000000110000011" => rgb <= "101111";
					when "000000110000100" => rgb <= "101111";
					when "000000110000101" => rgb <= "101111";
					when "000000110000110" => rgb <= "101111";
					when "000000110000111" => rgb <= "101111";
					when "000000110001000" => rgb <= "101111";
					when "000000110001001" => rgb <= "101111";
					when "000000110001010" => rgb <= "101111";
					when "000000110001011" => rgb <= "101111";
					when "000000110001100" => rgb <= "101111";
					when "000000110001101" => rgb <= "101111";
					when "000000110001110" => rgb <= "101111";
					when "000000110001111" => rgb <= "101111";
					when "000000110010000" => rgb <= "101111";
					when "000000110010001" => rgb <= "101111";
					when "000000110010010" => rgb <= "101111";
					when "000000110010011" => rgb <= "101111";
					when "000000110010100" => rgb <= "101111";
					when "000000110010101" => rgb <= "101111";
					when "000000110010110" => rgb <= "101111";
					when "000000110010111" => rgb <= "101111";
					when "000000110011000" => rgb <= "101111";
					when "000000110011001" => rgb <= "101111";
					when "000000110011010" => rgb <= "101111";
					when "000000110011011" => rgb <= "101111";
					when "000000110011100" => rgb <= "101111";
					when "000000110011101" => rgb <= "101111";
					when "000000110011110" => rgb <= "101111";
					when "000000110011111" => rgb <= "101111";
					when "000001000000000" => rgb <= "101111";
					when "000001000000001" => rgb <= "101111";
					when "000001000000010" => rgb <= "101111";
					when "000001000000011" => rgb <= "101111";
					when "000001000000100" => rgb <= "101111";
					when "000001000000101" => rgb <= "101111";
					when "000001000000110" => rgb <= "101111";
					when "000001000000111" => rgb <= "101111";
					when "000001000001000" => rgb <= "101111";
					when "000001000001001" => rgb <= "101111";
					when "000001000001010" => rgb <= "101111";
					when "000001000001011" => rgb <= "101111";
					when "000001000001100" => rgb <= "101111";
					when "000001000001101" => rgb <= "101111";
					when "000001000001110" => rgb <= "101111";
					when "000001000001111" => rgb <= "101111";
					when "000001000010000" => rgb <= "000000";
					when "000001000010001" => rgb <= "000000";
					when "000001000010010" => rgb <= "000000";
					when "000001000010011" => rgb <= "000000";
					when "000001000010100" => rgb <= "000000";
					when "000001000010101" => rgb <= "000000";
					when "000001000010110" => rgb <= "000000";
					when "000001000010111" => rgb <= "000000";
					when "000001000011000" => rgb <= "000000";
					when "000001000011001" => rgb <= "000000";
					when "000001000011010" => rgb <= "000000";
					when "000001000011011" => rgb <= "000000";
					when "000001000011100" => rgb <= "000000";
					when "000001000011101" => rgb <= "000000";
					when "000001000011110" => rgb <= "101111";
					when "000001000011111" => rgb <= "101111";
					when "000001000100000" => rgb <= "101111";
					when "000001000100001" => rgb <= "101111";
					when "000001000100010" => rgb <= "101111";
					when "000001000100011" => rgb <= "101111";
					when "000001000100100" => rgb <= "101111";
					when "000001000100101" => rgb <= "101111";
					when "000001000100110" => rgb <= "101111";
					when "000001000100111" => rgb <= "101111";
					when "000001000101000" => rgb <= "101111";
					when "000001000101001" => rgb <= "101111";
					when "000001000101010" => rgb <= "101111";
					when "000001000101011" => rgb <= "101111";
					when "000001000101100" => rgb <= "101111";
					when "000001000101101" => rgb <= "101111";
					when "000001000101110" => rgb <= "101111";
					when "000001000101111" => rgb <= "101111";
					when "000001000110000" => rgb <= "101111";
					when "000001000110001" => rgb <= "101111";
					when "000001000110010" => rgb <= "101111";
					when "000001000110011" => rgb <= "101111";
					when "000001000110100" => rgb <= "101111";
					when "000001000110101" => rgb <= "101111";
					when "000001000110110" => rgb <= "101111";
					when "000001000110111" => rgb <= "101111";
					when "000001000111000" => rgb <= "101111";
					when "000001000111001" => rgb <= "101111";
					when "000001000111010" => rgb <= "101111";
					when "000001000111011" => rgb <= "101111";
					when "000001000111100" => rgb <= "101111";
					when "000001000111101" => rgb <= "101111";
					when "000001000111110" => rgb <= "101111";
					when "000001000111111" => rgb <= "101111";
					when "000001001000000" => rgb <= "101111";
					when "000001001000001" => rgb <= "101111";
					when "000001001000010" => rgb <= "101111";
					when "000001001000011" => rgb <= "101111";
					when "000001001000100" => rgb <= "101111";
					when "000001001000101" => rgb <= "101111";
					when "000001001000110" => rgb <= "101111";
					when "000001001000111" => rgb <= "101111";
					when "000001001001000" => rgb <= "101111";
					when "000001001001001" => rgb <= "101111";
					when "000001001001010" => rgb <= "101111";
					when "000001001001011" => rgb <= "101111";
					when "000001001001100" => rgb <= "101111";
					when "000001001001101" => rgb <= "101111";
					when "000001001001110" => rgb <= "101111";
					when "000001001001111" => rgb <= "101111";
					when "000001001010000" => rgb <= "101111";
					when "000001001010001" => rgb <= "101111";
					when "000001001010010" => rgb <= "101111";
					when "000001001010011" => rgb <= "101111";
					when "000001001010100" => rgb <= "101111";
					when "000001001010101" => rgb <= "101111";
					when "000001001010110" => rgb <= "101111";
					when "000001001010111" => rgb <= "101111";
					when "000001001011000" => rgb <= "101111";
					when "000001001011001" => rgb <= "101111";
					when "000001001011010" => rgb <= "101111";
					when "000001001011011" => rgb <= "101111";
					when "000001001011100" => rgb <= "101111";
					when "000001001011101" => rgb <= "101111";
					when "000001001011110" => rgb <= "101111";
					when "000001001011111" => rgb <= "101111";
					when "000001001100000" => rgb <= "101111";
					when "000001001100001" => rgb <= "101111";
					when "000001001100010" => rgb <= "101111";
					when "000001001100011" => rgb <= "101111";
					when "000001001100100" => rgb <= "101111";
					when "000001001100101" => rgb <= "101111";
					when "000001001100110" => rgb <= "101111";
					when "000001001100111" => rgb <= "101111";
					when "000001001101000" => rgb <= "101111";
					when "000001001101001" => rgb <= "101111";
					when "000001001101010" => rgb <= "101111";
					when "000001001101011" => rgb <= "101111";
					when "000001001101100" => rgb <= "101111";
					when "000001001101101" => rgb <= "101111";
					when "000001001101110" => rgb <= "101111";
					when "000001001101111" => rgb <= "101111";
					when "000001001110000" => rgb <= "101111";
					when "000001001110001" => rgb <= "101111";
					when "000001001110010" => rgb <= "101111";
					when "000001001110011" => rgb <= "101111";
					when "000001001110100" => rgb <= "101111";
					when "000001001110101" => rgb <= "101111";
					when "000001001110110" => rgb <= "101111";
					when "000001001110111" => rgb <= "101111";
					when "000001001111000" => rgb <= "101111";
					when "000001001111001" => rgb <= "101111";
					when "000001001111010" => rgb <= "101111";
					when "000001001111011" => rgb <= "101111";
					when "000001001111100" => rgb <= "101111";
					when "000001001111101" => rgb <= "101111";
					when "000001001111110" => rgb <= "101111";
					when "000001001111111" => rgb <= "101111";
					when "000001010000000" => rgb <= "101111";
					when "000001010000001" => rgb <= "101111";
					when "000001010000010" => rgb <= "101111";
					when "000001010000011" => rgb <= "101111";
					when "000001010000100" => rgb <= "101111";
					when "000001010000101" => rgb <= "101111";
					when "000001010000110" => rgb <= "101111";
					when "000001010000111" => rgb <= "101111";
					when "000001010001000" => rgb <= "101111";
					when "000001010001001" => rgb <= "101111";
					when "000001010001010" => rgb <= "101111";
					when "000001010001011" => rgb <= "101111";
					when "000001010001100" => rgb <= "101111";
					when "000001010001101" => rgb <= "101111";
					when "000001010001110" => rgb <= "101111";
					when "000001010001111" => rgb <= "101111";
					when "000001010010000" => rgb <= "101111";
					when "000001010010001" => rgb <= "101111";
					when "000001010010010" => rgb <= "101111";
					when "000001010010011" => rgb <= "101111";
					when "000001010010100" => rgb <= "101111";
					when "000001010010101" => rgb <= "101111";
					when "000001010010110" => rgb <= "101111";
					when "000001010010111" => rgb <= "101111";
					when "000001010011000" => rgb <= "101111";
					when "000001010011001" => rgb <= "101111";
					when "000001010011010" => rgb <= "101111";
					when "000001010011011" => rgb <= "101111";
					when "000001010011100" => rgb <= "101111";
					when "000001010011101" => rgb <= "101111";
					when "000001010011110" => rgb <= "101111";
					when "000001010011111" => rgb <= "101111";
					when "000001100000000" => rgb <= "101111";
					when "000001100000001" => rgb <= "101111";
					when "000001100000010" => rgb <= "101111";
					when "000001100000011" => rgb <= "101111";
					when "000001100000100" => rgb <= "101111";
					when "000001100000101" => rgb <= "101111";
					when "000001100000110" => rgb <= "101111";
					when "000001100000111" => rgb <= "101111";
					when "000001100001000" => rgb <= "101111";
					when "000001100001001" => rgb <= "101111";
					when "000001100001010" => rgb <= "101111";
					when "000001100001011" => rgb <= "101111";
					when "000001100001100" => rgb <= "101111";
					when "000001100001101" => rgb <= "101111";
					when "000001100001110" => rgb <= "101111";
					when "000001100001111" => rgb <= "101111";
					when "000001100010000" => rgb <= "000000";
					when "000001100010001" => rgb <= "000000";
					when "000001100010010" => rgb <= "000000";
					when "000001100010011" => rgb <= "000000";
					when "000001100010100" => rgb <= "000000";
					when "000001100010101" => rgb <= "000000";
					when "000001100010110" => rgb <= "000000";
					when "000001100010111" => rgb <= "000000";
					when "000001100011000" => rgb <= "000000";
					when "000001100011001" => rgb <= "000000";
					when "000001100011010" => rgb <= "000000";
					when "000001100011011" => rgb <= "000000";
					when "000001100011100" => rgb <= "000000";
					when "000001100011101" => rgb <= "000000";
					when "000001100011110" => rgb <= "101111";
					when "000001100011111" => rgb <= "101111";
					when "000001100100000" => rgb <= "101111";
					when "000001100100001" => rgb <= "101111";
					when "000001100100010" => rgb <= "101111";
					when "000001100100011" => rgb <= "101111";
					when "000001100100100" => rgb <= "101111";
					when "000001100100101" => rgb <= "101111";
					when "000001100100110" => rgb <= "101111";
					when "000001100100111" => rgb <= "101111";
					when "000001100101000" => rgb <= "101111";
					when "000001100101001" => rgb <= "101111";
					when "000001100101010" => rgb <= "101111";
					when "000001100101011" => rgb <= "101111";
					when "000001100101100" => rgb <= "101111";
					when "000001100101101" => rgb <= "101111";
					when "000001100101110" => rgb <= "101111";
					when "000001100101111" => rgb <= "101111";
					when "000001100110000" => rgb <= "101111";
					when "000001100110001" => rgb <= "101111";
					when "000001100110010" => rgb <= "101111";
					when "000001100110011" => rgb <= "101111";
					when "000001100110100" => rgb <= "101111";
					when "000001100110101" => rgb <= "101111";
					when "000001100110110" => rgb <= "101111";
					when "000001100110111" => rgb <= "101111";
					when "000001100111000" => rgb <= "101111";
					when "000001100111001" => rgb <= "101111";
					when "000001100111010" => rgb <= "101111";
					when "000001100111011" => rgb <= "101111";
					when "000001100111100" => rgb <= "101111";
					when "000001100111101" => rgb <= "101111";
					when "000001100111110" => rgb <= "101111";
					when "000001100111111" => rgb <= "101111";
					when "000001101000000" => rgb <= "101111";
					when "000001101000001" => rgb <= "101111";
					when "000001101000010" => rgb <= "101111";
					when "000001101000011" => rgb <= "101111";
					when "000001101000100" => rgb <= "101111";
					when "000001101000101" => rgb <= "101111";
					when "000001101000110" => rgb <= "101111";
					when "000001101000111" => rgb <= "101111";
					when "000001101001000" => rgb <= "101111";
					when "000001101001001" => rgb <= "101111";
					when "000001101001010" => rgb <= "101111";
					when "000001101001011" => rgb <= "101111";
					when "000001101001100" => rgb <= "101111";
					when "000001101001101" => rgb <= "101111";
					when "000001101001110" => rgb <= "101111";
					when "000001101001111" => rgb <= "101111";
					when "000001101010000" => rgb <= "101111";
					when "000001101010001" => rgb <= "101111";
					when "000001101010010" => rgb <= "101111";
					when "000001101010011" => rgb <= "101111";
					when "000001101010100" => rgb <= "101111";
					when "000001101010101" => rgb <= "101111";
					when "000001101010110" => rgb <= "101111";
					when "000001101010111" => rgb <= "101111";
					when "000001101011000" => rgb <= "101111";
					when "000001101011001" => rgb <= "101111";
					when "000001101011010" => rgb <= "101111";
					when "000001101011011" => rgb <= "101111";
					when "000001101011100" => rgb <= "101111";
					when "000001101011101" => rgb <= "101111";
					when "000001101011110" => rgb <= "101111";
					when "000001101011111" => rgb <= "101111";
					when "000001101100000" => rgb <= "101111";
					when "000001101100001" => rgb <= "101111";
					when "000001101100010" => rgb <= "101111";
					when "000001101100011" => rgb <= "101111";
					when "000001101100100" => rgb <= "101111";
					when "000001101100101" => rgb <= "101111";
					when "000001101100110" => rgb <= "101111";
					when "000001101100111" => rgb <= "101111";
					when "000001101101000" => rgb <= "101111";
					when "000001101101001" => rgb <= "101111";
					when "000001101101010" => rgb <= "101111";
					when "000001101101011" => rgb <= "101111";
					when "000001101101100" => rgb <= "101111";
					when "000001101101101" => rgb <= "101111";
					when "000001101101110" => rgb <= "101111";
					when "000001101101111" => rgb <= "101111";
					when "000001101110000" => rgb <= "101111";
					when "000001101110001" => rgb <= "101111";
					when "000001101110010" => rgb <= "101111";
					when "000001101110011" => rgb <= "101111";
					when "000001101110100" => rgb <= "101111";
					when "000001101110101" => rgb <= "101111";
					when "000001101110110" => rgb <= "101111";
					when "000001101110111" => rgb <= "101111";
					when "000001101111000" => rgb <= "101111";
					when "000001101111001" => rgb <= "101111";
					when "000001101111010" => rgb <= "101111";
					when "000001101111011" => rgb <= "101111";
					when "000001101111100" => rgb <= "101111";
					when "000001101111101" => rgb <= "101111";
					when "000001101111110" => rgb <= "101111";
					when "000001101111111" => rgb <= "101111";
					when "000001110000000" => rgb <= "101111";
					when "000001110000001" => rgb <= "101111";
					when "000001110000010" => rgb <= "101111";
					when "000001110000011" => rgb <= "101111";
					when "000001110000100" => rgb <= "101111";
					when "000001110000101" => rgb <= "101111";
					when "000001110000110" => rgb <= "101111";
					when "000001110000111" => rgb <= "101111";
					when "000001110001000" => rgb <= "101111";
					when "000001110001001" => rgb <= "101111";
					when "000001110001010" => rgb <= "101111";
					when "000001110001011" => rgb <= "101111";
					when "000001110001100" => rgb <= "101111";
					when "000001110001101" => rgb <= "101111";
					when "000001110001110" => rgb <= "101111";
					when "000001110001111" => rgb <= "101111";
					when "000001110010000" => rgb <= "101111";
					when "000001110010001" => rgb <= "101111";
					when "000001110010010" => rgb <= "101111";
					when "000001110010011" => rgb <= "101111";
					when "000001110010100" => rgb <= "101111";
					when "000001110010101" => rgb <= "101111";
					when "000001110010110" => rgb <= "101111";
					when "000001110010111" => rgb <= "101111";
					when "000001110011000" => rgb <= "101111";
					when "000001110011001" => rgb <= "101111";
					when "000001110011010" => rgb <= "101111";
					when "000001110011011" => rgb <= "101111";
					when "000001110011100" => rgb <= "101111";
					when "000001110011101" => rgb <= "101111";
					when "000001110011110" => rgb <= "101111";
					when "000001110011111" => rgb <= "101111";
					when "000010000000000" => rgb <= "101111";
					when "000010000000001" => rgb <= "101111";
					when "000010000000010" => rgb <= "101111";
					when "000010000000011" => rgb <= "101111";
					when "000010000000100" => rgb <= "101111";
					when "000010000000101" => rgb <= "101111";
					when "000010000000110" => rgb <= "101111";
					when "000010000000111" => rgb <= "101111";
					when "000010000001000" => rgb <= "101111";
					when "000010000001001" => rgb <= "101111";
					when "000010000001010" => rgb <= "101111";
					when "000010000001011" => rgb <= "101111";
					when "000010000001100" => rgb <= "101111";
					when "000010000001101" => rgb <= "101111";
					when "000010000001110" => rgb <= "000000";
					when "000010000001111" => rgb <= "000000";
					when "000010000010000" => rgb <= "000000";
					when "000010000010001" => rgb <= "000000";
					when "000010000010010" => rgb <= "001000";
					when "000010000010011" => rgb <= "001000";
					when "000010000010100" => rgb <= "001000";
					when "000010000010101" => rgb <= "001000";
					when "000010000010110" => rgb <= "001000";
					when "000010000010111" => rgb <= "001000";
					when "000010000011000" => rgb <= "001000";
					when "000010000011001" => rgb <= "001000";
					when "000010000011010" => rgb <= "001000";
					when "000010000011011" => rgb <= "001000";
					when "000010000011100" => rgb <= "001000";
					when "000010000011101" => rgb <= "001000";
					when "000010000011110" => rgb <= "000000";
					when "000010000011111" => rgb <= "000000";
					when "000010000100000" => rgb <= "000000";
					when "000010000100001" => rgb <= "000000";
					when "000010000100010" => rgb <= "000000";
					when "000010000100011" => rgb <= "000000";
					when "000010000100100" => rgb <= "000000";
					when "000010000100101" => rgb <= "000000";
					when "000010000100110" => rgb <= "101111";
					when "000010000100111" => rgb <= "101111";
					when "000010000101000" => rgb <= "101111";
					when "000010000101001" => rgb <= "101111";
					when "000010000101010" => rgb <= "101111";
					when "000010000101011" => rgb <= "101111";
					when "000010000101100" => rgb <= "101111";
					when "000010000101101" => rgb <= "101111";
					when "000010000101110" => rgb <= "101111";
					when "000010000101111" => rgb <= "101111";
					when "000010000110000" => rgb <= "101111";
					when "000010000110001" => rgb <= "101111";
					when "000010000110010" => rgb <= "101111";
					when "000010000110011" => rgb <= "101111";
					when "000010000110100" => rgb <= "101111";
					when "000010000110101" => rgb <= "101111";
					when "000010000110110" => rgb <= "101111";
					when "000010000110111" => rgb <= "101111";
					when "000010000111000" => rgb <= "101111";
					when "000010000111001" => rgb <= "101111";
					when "000010000111010" => rgb <= "101111";
					when "000010000111011" => rgb <= "101111";
					when "000010000111100" => rgb <= "101111";
					when "000010000111101" => rgb <= "101111";
					when "000010000111110" => rgb <= "101111";
					when "000010000111111" => rgb <= "101111";
					when "000010001000000" => rgb <= "101111";
					when "000010001000001" => rgb <= "101111";
					when "000010001000010" => rgb <= "101111";
					when "000010001000011" => rgb <= "101111";
					when "000010001000100" => rgb <= "101111";
					when "000010001000101" => rgb <= "101111";
					when "000010001000110" => rgb <= "101111";
					when "000010001000111" => rgb <= "101111";
					when "000010001001000" => rgb <= "101111";
					when "000010001001001" => rgb <= "101111";
					when "000010001001010" => rgb <= "101111";
					when "000010001001011" => rgb <= "101111";
					when "000010001001100" => rgb <= "101111";
					when "000010001001101" => rgb <= "101111";
					when "000010001001110" => rgb <= "101111";
					when "000010001001111" => rgb <= "101111";
					when "000010001010000" => rgb <= "101111";
					when "000010001010001" => rgb <= "101111";
					when "000010001010010" => rgb <= "101111";
					when "000010001010011" => rgb <= "101111";
					when "000010001010100" => rgb <= "101111";
					when "000010001010101" => rgb <= "101111";
					when "000010001010110" => rgb <= "101111";
					when "000010001010111" => rgb <= "101111";
					when "000010001011000" => rgb <= "101111";
					when "000010001011001" => rgb <= "101111";
					when "000010001011010" => rgb <= "101111";
					when "000010001011011" => rgb <= "101111";
					when "000010001011100" => rgb <= "101111";
					when "000010001011101" => rgb <= "101111";
					when "000010001011110" => rgb <= "101111";
					when "000010001011111" => rgb <= "101111";
					when "000010001100000" => rgb <= "101111";
					when "000010001100001" => rgb <= "101111";
					when "000010001100010" => rgb <= "101111";
					when "000010001100011" => rgb <= "101111";
					when "000010001100100" => rgb <= "101111";
					when "000010001100101" => rgb <= "101111";
					when "000010001100110" => rgb <= "101111";
					when "000010001100111" => rgb <= "101111";
					when "000010001101000" => rgb <= "101111";
					when "000010001101001" => rgb <= "101111";
					when "000010001101010" => rgb <= "101111";
					when "000010001101011" => rgb <= "101111";
					when "000010001101100" => rgb <= "101111";
					when "000010001101101" => rgb <= "101111";
					when "000010001101110" => rgb <= "101111";
					when "000010001101111" => rgb <= "101111";
					when "000010001110000" => rgb <= "101111";
					when "000010001110001" => rgb <= "101111";
					when "000010001110010" => rgb <= "101111";
					when "000010001110011" => rgb <= "101111";
					when "000010001110100" => rgb <= "101111";
					when "000010001110101" => rgb <= "101111";
					when "000010001110110" => rgb <= "101111";
					when "000010001110111" => rgb <= "101111";
					when "000010001111000" => rgb <= "101111";
					when "000010001111001" => rgb <= "101111";
					when "000010001111010" => rgb <= "101111";
					when "000010001111011" => rgb <= "101111";
					when "000010001111100" => rgb <= "101111";
					when "000010001111101" => rgb <= "101111";
					when "000010001111110" => rgb <= "101111";
					when "000010001111111" => rgb <= "101111";
					when "000010010000000" => rgb <= "101111";
					when "000010010000001" => rgb <= "101111";
					when "000010010000010" => rgb <= "101111";
					when "000010010000011" => rgb <= "101111";
					when "000010010000100" => rgb <= "101111";
					when "000010010000101" => rgb <= "101111";
					when "000010010000110" => rgb <= "101111";
					when "000010010000111" => rgb <= "101111";
					when "000010010001000" => rgb <= "101111";
					when "000010010001001" => rgb <= "101111";
					when "000010010001010" => rgb <= "101111";
					when "000010010001011" => rgb <= "101111";
					when "000010010001100" => rgb <= "101111";
					when "000010010001101" => rgb <= "101111";
					when "000010010001110" => rgb <= "101111";
					when "000010010001111" => rgb <= "101111";
					when "000010010010000" => rgb <= "101111";
					when "000010010010001" => rgb <= "101111";
					when "000010010010010" => rgb <= "101111";
					when "000010010010011" => rgb <= "101111";
					when "000010010010100" => rgb <= "101111";
					when "000010010010101" => rgb <= "101111";
					when "000010010010110" => rgb <= "101111";
					when "000010010010111" => rgb <= "101111";
					when "000010010011000" => rgb <= "101111";
					when "000010010011001" => rgb <= "101111";
					when "000010010011010" => rgb <= "101111";
					when "000010010011011" => rgb <= "101111";
					when "000010010011100" => rgb <= "101111";
					when "000010010011101" => rgb <= "101111";
					when "000010010011110" => rgb <= "101111";
					when "000010010011111" => rgb <= "101111";
					when "000010100000000" => rgb <= "101111";
					when "000010100000001" => rgb <= "101111";
					when "000010100000010" => rgb <= "101111";
					when "000010100000011" => rgb <= "101111";
					when "000010100000100" => rgb <= "101111";
					when "000010100000101" => rgb <= "101111";
					when "000010100000110" => rgb <= "101111";
					when "000010100000111" => rgb <= "101111";
					when "000010100001000" => rgb <= "101111";
					when "000010100001001" => rgb <= "101111";
					when "000010100001010" => rgb <= "101111";
					when "000010100001011" => rgb <= "101111";
					when "000010100001100" => rgb <= "101111";
					when "000010100001101" => rgb <= "101111";
					when "000010100001110" => rgb <= "000000";
					when "000010100001111" => rgb <= "000000";
					when "000010100010000" => rgb <= "000000";
					when "000010100010001" => rgb <= "000000";
					when "000010100010010" => rgb <= "001000";
					when "000010100010011" => rgb <= "001000";
					when "000010100010100" => rgb <= "001000";
					when "000010100010101" => rgb <= "001000";
					when "000010100010110" => rgb <= "001000";
					when "000010100010111" => rgb <= "001000";
					when "000010100011000" => rgb <= "001000";
					when "000010100011001" => rgb <= "001000";
					when "000010100011010" => rgb <= "001000";
					when "000010100011011" => rgb <= "001000";
					when "000010100011100" => rgb <= "001000";
					when "000010100011101" => rgb <= "001000";
					when "000010100011110" => rgb <= "000000";
					when "000010100011111" => rgb <= "000000";
					when "000010100100000" => rgb <= "000000";
					when "000010100100001" => rgb <= "000000";
					when "000010100100010" => rgb <= "000000";
					when "000010100100011" => rgb <= "000000";
					when "000010100100100" => rgb <= "000000";
					when "000010100100101" => rgb <= "000000";
					when "000010100100110" => rgb <= "101111";
					when "000010100100111" => rgb <= "101111";
					when "000010100101000" => rgb <= "101111";
					when "000010100101001" => rgb <= "101111";
					when "000010100101010" => rgb <= "101111";
					when "000010100101011" => rgb <= "101111";
					when "000010100101100" => rgb <= "101111";
					when "000010100101101" => rgb <= "101111";
					when "000010100101110" => rgb <= "101111";
					when "000010100101111" => rgb <= "101111";
					when "000010100110000" => rgb <= "101111";
					when "000010100110001" => rgb <= "101111";
					when "000010100110010" => rgb <= "101111";
					when "000010100110011" => rgb <= "101111";
					when "000010100110100" => rgb <= "101111";
					when "000010100110101" => rgb <= "101111";
					when "000010100110110" => rgb <= "101111";
					when "000010100110111" => rgb <= "101111";
					when "000010100111000" => rgb <= "101111";
					when "000010100111001" => rgb <= "101111";
					when "000010100111010" => rgb <= "101111";
					when "000010100111011" => rgb <= "101111";
					when "000010100111100" => rgb <= "101111";
					when "000010100111101" => rgb <= "101111";
					when "000010100111110" => rgb <= "101111";
					when "000010100111111" => rgb <= "101111";
					when "000010101000000" => rgb <= "101111";
					when "000010101000001" => rgb <= "101111";
					when "000010101000010" => rgb <= "101111";
					when "000010101000011" => rgb <= "101111";
					when "000010101000100" => rgb <= "101111";
					when "000010101000101" => rgb <= "101111";
					when "000010101000110" => rgb <= "101111";
					when "000010101000111" => rgb <= "101111";
					when "000010101001000" => rgb <= "101111";
					when "000010101001001" => rgb <= "101111";
					when "000010101001010" => rgb <= "101111";
					when "000010101001011" => rgb <= "101111";
					when "000010101001100" => rgb <= "101111";
					when "000010101001101" => rgb <= "101111";
					when "000010101001110" => rgb <= "101111";
					when "000010101001111" => rgb <= "101111";
					when "000010101010000" => rgb <= "101111";
					when "000010101010001" => rgb <= "101111";
					when "000010101010010" => rgb <= "101111";
					when "000010101010011" => rgb <= "101111";
					when "000010101010100" => rgb <= "101111";
					when "000010101010101" => rgb <= "101111";
					when "000010101010110" => rgb <= "101111";
					when "000010101010111" => rgb <= "101111";
					when "000010101011000" => rgb <= "101111";
					when "000010101011001" => rgb <= "101111";
					when "000010101011010" => rgb <= "101111";
					when "000010101011011" => rgb <= "101111";
					when "000010101011100" => rgb <= "101111";
					when "000010101011101" => rgb <= "101111";
					when "000010101011110" => rgb <= "101111";
					when "000010101011111" => rgb <= "101111";
					when "000010101100000" => rgb <= "101111";
					when "000010101100001" => rgb <= "101111";
					when "000010101100010" => rgb <= "101111";
					when "000010101100011" => rgb <= "101111";
					when "000010101100100" => rgb <= "101111";
					when "000010101100101" => rgb <= "101111";
					when "000010101100110" => rgb <= "101111";
					when "000010101100111" => rgb <= "101111";
					when "000010101101000" => rgb <= "101111";
					when "000010101101001" => rgb <= "101111";
					when "000010101101010" => rgb <= "101111";
					when "000010101101011" => rgb <= "101111";
					when "000010101101100" => rgb <= "101111";
					when "000010101101101" => rgb <= "101111";
					when "000010101101110" => rgb <= "101111";
					when "000010101101111" => rgb <= "101111";
					when "000010101110000" => rgb <= "101111";
					when "000010101110001" => rgb <= "101111";
					when "000010101110010" => rgb <= "101111";
					when "000010101110011" => rgb <= "101111";
					when "000010101110100" => rgb <= "101111";
					when "000010101110101" => rgb <= "101111";
					when "000010101110110" => rgb <= "101111";
					when "000010101110111" => rgb <= "101111";
					when "000010101111000" => rgb <= "101111";
					when "000010101111001" => rgb <= "101111";
					when "000010101111010" => rgb <= "101111";
					when "000010101111011" => rgb <= "101111";
					when "000010101111100" => rgb <= "101111";
					when "000010101111101" => rgb <= "101111";
					when "000010101111110" => rgb <= "101111";
					when "000010101111111" => rgb <= "101111";
					when "000010110000000" => rgb <= "101111";
					when "000010110000001" => rgb <= "101111";
					when "000010110000010" => rgb <= "101111";
					when "000010110000011" => rgb <= "101111";
					when "000010110000100" => rgb <= "101111";
					when "000010110000101" => rgb <= "101111";
					when "000010110000110" => rgb <= "101111";
					when "000010110000111" => rgb <= "101111";
					when "000010110001000" => rgb <= "101111";
					when "000010110001001" => rgb <= "101111";
					when "000010110001010" => rgb <= "101111";
					when "000010110001011" => rgb <= "101111";
					when "000010110001100" => rgb <= "101111";
					when "000010110001101" => rgb <= "101111";
					when "000010110001110" => rgb <= "101111";
					when "000010110001111" => rgb <= "101111";
					when "000010110010000" => rgb <= "101111";
					when "000010110010001" => rgb <= "101111";
					when "000010110010010" => rgb <= "101111";
					when "000010110010011" => rgb <= "101111";
					when "000010110010100" => rgb <= "101111";
					when "000010110010101" => rgb <= "101111";
					when "000010110010110" => rgb <= "101111";
					when "000010110010111" => rgb <= "101111";
					when "000010110011000" => rgb <= "101111";
					when "000010110011001" => rgb <= "101111";
					when "000010110011010" => rgb <= "101111";
					when "000010110011011" => rgb <= "101111";
					when "000010110011100" => rgb <= "101111";
					when "000010110011101" => rgb <= "101111";
					when "000010110011110" => rgb <= "101111";
					when "000010110011111" => rgb <= "101111";
					when "000011000000000" => rgb <= "101111";
					when "000011000000001" => rgb <= "101111";
					when "000011000000010" => rgb <= "101111";
					when "000011000000011" => rgb <= "101111";
					when "000011000000100" => rgb <= "101111";
					when "000011000000101" => rgb <= "101111";
					when "000011000000110" => rgb <= "101111";
					when "000011000000111" => rgb <= "101111";
					when "000011000001000" => rgb <= "101111";
					when "000011000001001" => rgb <= "101111";
					when "000011000001010" => rgb <= "101111";
					when "000011000001011" => rgb <= "101111";
					when "000011000001100" => rgb <= "101111";
					when "000011000001101" => rgb <= "101111";
					when "000011000001110" => rgb <= "101111";
					when "000011000001111" => rgb <= "000000";
					when "000011000010000" => rgb <= "101111";
					when "000011000010001" => rgb <= "101111";
					when "000011000010010" => rgb <= "101111";
					when "000011000010011" => rgb <= "101111";
					when "000011000010100" => rgb <= "101111";
					when "000011000010101" => rgb <= "001000";
					when "000011000010110" => rgb <= "001000";
					when "000011000010111" => rgb <= "101111";
					when "000011000011000" => rgb <= "101111";
					when "000011000011001" => rgb <= "101111";
					when "000011000011010" => rgb <= "101111";
					when "000011000011011" => rgb <= "101111";
					when "000011000011100" => rgb <= "101111";
					when "000011000011101" => rgb <= "101111";
					when "000011000011110" => rgb <= "001000";
					when "000011000011111" => rgb <= "101111";
					when "000011000100000" => rgb <= "101111";
					when "000011000100001" => rgb <= "101111";
					when "000011000100010" => rgb <= "101111";
					when "000011000100011" => rgb <= "101111";
					when "000011000100100" => rgb <= "101111";
					when "000011000100101" => rgb <= "101111";
					when "000011000100110" => rgb <= "101111";
					when "000011000100111" => rgb <= "101111";
					when "000011000101000" => rgb <= "000000";
					when "000011000101001" => rgb <= "000000";
					when "000011000101010" => rgb <= "000000";
					when "000011000101011" => rgb <= "000000";
					when "000011000101100" => rgb <= "000000";
					when "000011000101101" => rgb <= "000000";
					when "000011000101110" => rgb <= "000000";
					when "000011000101111" => rgb <= "000000";
					when "000011000110000" => rgb <= "000000";
					when "000011000110001" => rgb <= "000000";
					when "000011000110010" => rgb <= "000000";
					when "000011000110011" => rgb <= "000000";
					when "000011000110100" => rgb <= "000000";
					when "000011000110101" => rgb <= "000000";
					when "000011000110110" => rgb <= "000000";
					when "000011000110111" => rgb <= "000000";
					when "000011000111000" => rgb <= "000000";
					when "000011000111001" => rgb <= "000000";
					when "000011000111010" => rgb <= "000000";
					when "000011000111011" => rgb <= "000000";
					when "000011000111100" => rgb <= "000000";
					when "000011000111101" => rgb <= "000000";
					when "000011000111110" => rgb <= "000000";
					when "000011000111111" => rgb <= "000000";
					when "000011001000000" => rgb <= "000000";
					when "000011001000001" => rgb <= "000000";
					when "000011001000010" => rgb <= "000000";
					when "000011001000011" => rgb <= "000000";
					when "000011001000100" => rgb <= "000000";
					when "000011001000101" => rgb <= "000000";
					when "000011001000110" => rgb <= "000000";
					when "000011001000111" => rgb <= "000000";
					when "000011001001000" => rgb <= "000000";
					when "000011001001001" => rgb <= "000000";
					when "000011001001010" => rgb <= "000000";
					when "000011001001011" => rgb <= "000000";
					when "000011001001100" => rgb <= "000000";
					when "000011001001101" => rgb <= "000000";
					when "000011001001110" => rgb <= "000000";
					when "000011001001111" => rgb <= "000000";
					when "000011001010000" => rgb <= "000000";
					when "000011001010001" => rgb <= "000000";
					when "000011001010010" => rgb <= "000000";
					when "000011001010011" => rgb <= "000000";
					when "000011001010100" => rgb <= "000000";
					when "000011001010101" => rgb <= "000000";
					when "000011001010110" => rgb <= "000000";
					when "000011001010111" => rgb <= "000000";
					when "000011001011000" => rgb <= "000000";
					when "000011001011001" => rgb <= "000000";
					when "000011001011010" => rgb <= "000000";
					when "000011001011011" => rgb <= "000000";
					when "000011001011100" => rgb <= "000000";
					when "000011001011101" => rgb <= "000000";
					when "000011001011110" => rgb <= "000000";
					when "000011001011111" => rgb <= "000000";
					when "000011001100000" => rgb <= "000000";
					when "000011001100001" => rgb <= "000000";
					when "000011001100010" => rgb <= "000000";
					when "000011001100011" => rgb <= "000000";
					when "000011001100100" => rgb <= "000000";
					when "000011001100101" => rgb <= "000000";
					when "000011001100110" => rgb <= "000000";
					when "000011001100111" => rgb <= "000000";
					when "000011001101000" => rgb <= "000000";
					when "000011001101001" => rgb <= "000000";
					when "000011001101010" => rgb <= "000000";
					when "000011001101011" => rgb <= "000000";
					when "000011001101100" => rgb <= "000000";
					when "000011001101101" => rgb <= "000000";
					when "000011001101110" => rgb <= "000000";
					when "000011001101111" => rgb <= "000000";
					when "000011001110000" => rgb <= "000000";
					when "000011001110001" => rgb <= "000000";
					when "000011001110010" => rgb <= "000000";
					when "000011001110011" => rgb <= "000000";
					when "000011001110100" => rgb <= "000000";
					when "000011001110101" => rgb <= "000000";
					when "000011001110110" => rgb <= "000000";
					when "000011001110111" => rgb <= "000000";
					when "000011001111000" => rgb <= "101111";
					when "000011001111001" => rgb <= "101111";
					when "000011001111010" => rgb <= "101111";
					when "000011001111011" => rgb <= "101111";
					when "000011001111100" => rgb <= "101111";
					when "000011001111101" => rgb <= "101111";
					when "000011001111110" => rgb <= "101111";
					when "000011001111111" => rgb <= "101111";
					when "000011010000000" => rgb <= "101111";
					when "000011010000001" => rgb <= "101111";
					when "000011010000010" => rgb <= "101111";
					when "000011010000011" => rgb <= "101111";
					when "000011010000100" => rgb <= "101111";
					when "000011010000101" => rgb <= "101111";
					when "000011010000110" => rgb <= "101111";
					when "000011010000111" => rgb <= "101111";
					when "000011010001000" => rgb <= "101111";
					when "000011010001001" => rgb <= "101111";
					when "000011010001010" => rgb <= "101111";
					when "000011010001011" => rgb <= "101111";
					when "000011010001100" => rgb <= "101111";
					when "000011010001101" => rgb <= "101111";
					when "000011010001110" => rgb <= "101111";
					when "000011010001111" => rgb <= "101111";
					when "000011010010000" => rgb <= "101111";
					when "000011010010001" => rgb <= "101111";
					when "000011010010010" => rgb <= "101111";
					when "000011010010011" => rgb <= "101111";
					when "000011010010100" => rgb <= "101111";
					when "000011010010101" => rgb <= "101111";
					when "000011010010110" => rgb <= "101111";
					when "000011010010111" => rgb <= "101111";
					when "000011010011000" => rgb <= "101111";
					when "000011010011001" => rgb <= "101111";
					when "000011010011010" => rgb <= "101111";
					when "000011010011011" => rgb <= "101111";
					when "000011010011100" => rgb <= "101111";
					when "000011010011101" => rgb <= "101111";
					when "000011010011110" => rgb <= "101111";
					when "000011010011111" => rgb <= "101111";
					when "000011100000000" => rgb <= "101111";
					when "000011100000001" => rgb <= "101111";
					when "000011100000010" => rgb <= "101111";
					when "000011100000011" => rgb <= "101111";
					when "000011100000100" => rgb <= "101111";
					when "000011100000101" => rgb <= "101111";
					when "000011100000110" => rgb <= "101111";
					when "000011100000111" => rgb <= "000000";
					when "000011100001000" => rgb <= "000000";
					when "000011100001001" => rgb <= "000000";
					when "000011100001010" => rgb <= "000000";
					when "000011100001011" => rgb <= "000000";
					when "000011100001100" => rgb <= "000000";
					when "000011100001101" => rgb <= "101111";
					when "000011100001110" => rgb <= "101111";
					when "000011100001111" => rgb <= "101111";
					when "000011100010000" => rgb <= "101111";
					when "000011100010001" => rgb <= "000000";
					when "000011100010010" => rgb <= "000000";
					when "000011100010011" => rgb <= "000000";
					when "000011100010100" => rgb <= "101111";
					when "000011100010101" => rgb <= "101111";
					when "000011100010110" => rgb <= "001000";
					when "000011100010111" => rgb <= "101111";
					when "000011100011000" => rgb <= "000000";
					when "000011100011001" => rgb <= "101111";
					when "000011100011010" => rgb <= "101111";
					when "000011100011011" => rgb <= "000000";
					when "000011100011100" => rgb <= "000000";
					when "000011100011101" => rgb <= "101111";
					when "000011100011110" => rgb <= "101111";
					when "000011100011111" => rgb <= "101111";
					when "000011100100000" => rgb <= "000000";
					when "000011100100001" => rgb <= "000000";
					when "000011100100010" => rgb <= "101111";
					when "000011100100011" => rgb <= "101111";
					when "000011100100100" => rgb <= "000000";
					when "000011100100101" => rgb <= "000000";
					when "000011100100110" => rgb <= "000000";
					when "000011100100111" => rgb <= "101111";
					when "000011100101000" => rgb <= "000000";
					when "000011100101001" => rgb <= "000000";
					when "000011100101010" => rgb <= "000000";
					when "000011100101011" => rgb <= "000000";
					when "000011100101100" => rgb <= "000000";
					when "000011100101101" => rgb <= "000000";
					when "000011100101110" => rgb <= "000000";
					when "000011100101111" => rgb <= "000000";
					when "000011100110000" => rgb <= "000000";
					when "000011100110001" => rgb <= "000000";
					when "000011100110010" => rgb <= "000000";
					when "000011100110011" => rgb <= "000000";
					when "000011100110100" => rgb <= "000000";
					when "000011100110101" => rgb <= "000000";
					when "000011100110110" => rgb <= "000000";
					when "000011100110111" => rgb <= "000000";
					when "000011100111000" => rgb <= "000000";
					when "000011100111001" => rgb <= "000000";
					when "000011100111010" => rgb <= "000000";
					when "000011100111011" => rgb <= "000000";
					when "000011100111100" => rgb <= "000000";
					when "000011100111101" => rgb <= "000000";
					when "000011100111110" => rgb <= "000000";
					when "000011100111111" => rgb <= "000000";
					when "000011101000000" => rgb <= "000000";
					when "000011101000001" => rgb <= "000000";
					when "000011101000010" => rgb <= "000000";
					when "000011101000011" => rgb <= "000000";
					when "000011101000100" => rgb <= "000000";
					when "000011101000101" => rgb <= "000000";
					when "000011101000110" => rgb <= "000000";
					when "000011101000111" => rgb <= "000000";
					when "000011101001000" => rgb <= "000000";
					when "000011101001001" => rgb <= "000000";
					when "000011101001010" => rgb <= "000000";
					when "000011101001011" => rgb <= "000000";
					when "000011101001100" => rgb <= "000000";
					when "000011101001101" => rgb <= "000000";
					when "000011101001110" => rgb <= "000000";
					when "000011101001111" => rgb <= "000000";
					when "000011101010000" => rgb <= "000000";
					when "000011101010001" => rgb <= "000000";
					when "000011101010010" => rgb <= "000000";
					when "000011101010011" => rgb <= "000000";
					when "000011101010100" => rgb <= "000000";
					when "000011101010101" => rgb <= "000000";
					when "000011101010110" => rgb <= "000000";
					when "000011101010111" => rgb <= "000000";
					when "000011101011000" => rgb <= "000000";
					when "000011101011001" => rgb <= "000000";
					when "000011101011010" => rgb <= "000000";
					when "000011101011011" => rgb <= "000000";
					when "000011101011100" => rgb <= "000000";
					when "000011101011101" => rgb <= "000000";
					when "000011101011110" => rgb <= "000000";
					when "000011101011111" => rgb <= "000000";
					when "000011101100000" => rgb <= "000000";
					when "000011101100001" => rgb <= "000000";
					when "000011101100010" => rgb <= "000000";
					when "000011101100011" => rgb <= "000000";
					when "000011101100100" => rgb <= "000000";
					when "000011101100101" => rgb <= "000000";
					when "000011101100110" => rgb <= "000000";
					when "000011101100111" => rgb <= "000000";
					when "000011101101000" => rgb <= "000000";
					when "000011101101001" => rgb <= "000000";
					when "000011101101010" => rgb <= "000000";
					when "000011101101011" => rgb <= "000000";
					when "000011101101100" => rgb <= "000000";
					when "000011101101101" => rgb <= "000000";
					when "000011101101110" => rgb <= "000000";
					when "000011101101111" => rgb <= "000000";
					when "000011101110000" => rgb <= "000000";
					when "000011101110001" => rgb <= "000000";
					when "000011101110010" => rgb <= "000000";
					when "000011101110011" => rgb <= "000000";
					when "000011101110100" => rgb <= "000000";
					when "000011101110101" => rgb <= "000000";
					when "000011101110110" => rgb <= "000000";
					when "000011101110111" => rgb <= "000000";
					when "000011101111000" => rgb <= "101111";
					when "000011101111001" => rgb <= "101111";
					when "000011101111010" => rgb <= "000000";
					when "000011101111011" => rgb <= "000000";
					when "000011101111100" => rgb <= "000000";
					when "000011101111101" => rgb <= "000000";
					when "000011101111110" => rgb <= "000000";
					when "000011101111111" => rgb <= "101111";
					when "000011110000000" => rgb <= "101111";
					when "000011110000001" => rgb <= "101111";
					when "000011110000010" => rgb <= "000000";
					when "000011110000011" => rgb <= "000000";
					when "000011110000100" => rgb <= "101111";
					when "000011110000101" => rgb <= "101111";
					when "000011110000110" => rgb <= "000000";
					when "000011110000111" => rgb <= "000000";
					when "000011110001000" => rgb <= "101111";
					when "000011110001001" => rgb <= "101111";
					when "000011110001010" => rgb <= "101111";
					when "000011110001011" => rgb <= "000000";
					when "000011110001100" => rgb <= "101111";
					when "000011110001101" => rgb <= "101111";
					when "000011110001110" => rgb <= "000000";
					when "000011110001111" => rgb <= "000000";
					when "000011110010000" => rgb <= "101111";
					when "000011110010001" => rgb <= "101111";
					when "000011110010010" => rgb <= "101111";
					when "000011110010011" => rgb <= "000000";
					when "000011110010100" => rgb <= "000000";
					when "000011110010101" => rgb <= "000000";
					when "000011110010110" => rgb <= "000000";
					when "000011110010111" => rgb <= "101111";
					when "000011110011000" => rgb <= "101111";
					when "000011110011001" => rgb <= "101111";
					when "000011110011010" => rgb <= "000000";
					when "000011110011011" => rgb <= "000000";
					when "000011110011100" => rgb <= "101111";
					when "000011110011101" => rgb <= "101111";
					when "000011110011110" => rgb <= "101111";
					when "000011110011111" => rgb <= "101111";
					when "000100000000000" => rgb <= "101111";
					when "000100000000001" => rgb <= "101111";
					when "000100000000010" => rgb <= "101111";
					when "000100000000011" => rgb <= "101111";
					when "000100000000100" => rgb <= "101111";
					when "000100000000101" => rgb <= "101111";
					when "000100000000110" => rgb <= "000000";
					when "000100000000111" => rgb <= "110000";
					when "000100000001000" => rgb <= "110000";
					when "000100000001001" => rgb <= "110000";
					when "000100000001010" => rgb <= "110000";
					when "000100000001011" => rgb <= "110000";
					when "000100000001100" => rgb <= "110000";
					when "000100000001101" => rgb <= "000000";
					when "000100000001110" => rgb <= "101111";
					when "000100000001111" => rgb <= "101111";
					when "000100000010000" => rgb <= "000000";
					when "000100000010001" => rgb <= "110000";
					when "000100000010010" => rgb <= "110000";
					when "000100000010011" => rgb <= "110000";
					when "000100000010100" => rgb <= "000000";
					when "000100000010101" => rgb <= "101111";
					when "000100000010110" => rgb <= "101111";
					when "000100000010111" => rgb <= "000000";
					when "000100000011000" => rgb <= "110000";
					when "000100000011001" => rgb <= "000000";
					when "000100000011010" => rgb <= "000000";
					when "000100000011011" => rgb <= "110000";
					when "000100000011100" => rgb <= "110000";
					when "000100000011101" => rgb <= "000000";
					when "000100000011110" => rgb <= "101111";
					when "000100000011111" => rgb <= "000000";
					when "000100000100000" => rgb <= "110000";
					when "000100000100001" => rgb <= "110000";
					when "000100000100010" => rgb <= "000000";
					when "000100000100011" => rgb <= "000000";
					when "000100000100100" => rgb <= "110000";
					when "000100000100101" => rgb <= "110000";
					when "000100000100110" => rgb <= "000000";
					when "000100000100111" => rgb <= "101111";
					when "000100000101000" => rgb <= "000000";
					when "000100000101001" => rgb <= "000000";
					when "000100000101010" => rgb <= "101111";
					when "000100000101011" => rgb <= "101111";
					when "000100000101100" => rgb <= "101111";
					when "000100000101101" => rgb <= "101111";
					when "000100000101110" => rgb <= "101111";
					when "000100000101111" => rgb <= "101111";
					when "000100000110000" => rgb <= "101111";
					when "000100000110001" => rgb <= "101111";
					when "000100000110010" => rgb <= "101111";
					when "000100000110011" => rgb <= "101111";
					when "000100000110100" => rgb <= "101111";
					when "000100000110101" => rgb <= "101111";
					when "000100000110110" => rgb <= "101111";
					when "000100000110111" => rgb <= "101111";
					when "000100000111000" => rgb <= "101111";
					when "000100000111001" => rgb <= "101111";
					when "000100000111010" => rgb <= "101111";
					when "000100000111011" => rgb <= "101111";
					when "000100000111100" => rgb <= "101111";
					when "000100000111101" => rgb <= "101111";
					when "000100000111110" => rgb <= "101111";
					when "000100000111111" => rgb <= "101111";
					when "000100001000000" => rgb <= "101111";
					when "000100001000001" => rgb <= "101111";
					when "000100001000010" => rgb <= "101111";
					when "000100001000011" => rgb <= "101111";
					when "000100001000100" => rgb <= "101111";
					when "000100001000101" => rgb <= "101111";
					when "000100001000110" => rgb <= "101111";
					when "000100001000111" => rgb <= "101111";
					when "000100001001000" => rgb <= "101111";
					when "000100001001001" => rgb <= "101111";
					when "000100001001010" => rgb <= "101111";
					when "000100001001011" => rgb <= "101111";
					when "000100001001100" => rgb <= "101111";
					when "000100001001101" => rgb <= "101111";
					when "000100001001110" => rgb <= "101111";
					when "000100001001111" => rgb <= "101111";
					when "000100001010000" => rgb <= "101111";
					when "000100001010001" => rgb <= "101111";
					when "000100001010010" => rgb <= "101111";
					when "000100001010011" => rgb <= "101111";
					when "000100001010100" => rgb <= "101111";
					when "000100001010101" => rgb <= "101111";
					when "000100001010110" => rgb <= "101111";
					when "000100001010111" => rgb <= "101111";
					when "000100001011000" => rgb <= "101111";
					when "000100001011001" => rgb <= "101111";
					when "000100001011010" => rgb <= "101111";
					when "000100001011011" => rgb <= "101111";
					when "000100001011100" => rgb <= "101111";
					when "000100001011101" => rgb <= "101111";
					when "000100001011110" => rgb <= "101111";
					when "000100001011111" => rgb <= "101111";
					when "000100001100000" => rgb <= "101111";
					when "000100001100001" => rgb <= "101111";
					when "000100001100010" => rgb <= "101111";
					when "000100001100011" => rgb <= "101111";
					when "000100001100100" => rgb <= "101111";
					when "000100001100101" => rgb <= "101111";
					when "000100001100110" => rgb <= "101111";
					when "000100001100111" => rgb <= "101111";
					when "000100001101000" => rgb <= "101111";
					when "000100001101001" => rgb <= "101111";
					when "000100001101010" => rgb <= "101111";
					when "000100001101011" => rgb <= "101111";
					when "000100001101100" => rgb <= "101111";
					when "000100001101101" => rgb <= "101111";
					when "000100001101110" => rgb <= "101111";
					when "000100001101111" => rgb <= "101111";
					when "000100001110000" => rgb <= "101111";
					when "000100001110001" => rgb <= "101111";
					when "000100001110010" => rgb <= "101111";
					when "000100001110011" => rgb <= "101111";
					when "000100001110100" => rgb <= "101111";
					when "000100001110101" => rgb <= "101111";
					when "000100001110110" => rgb <= "000000";
					when "000100001110111" => rgb <= "000000";
					when "000100001111000" => rgb <= "101111";
					when "000100001111001" => rgb <= "000000";
					when "000100001111010" => rgb <= "000111";
					when "000100001111011" => rgb <= "000111";
					when "000100001111100" => rgb <= "000111";
					when "000100001111101" => rgb <= "000111";
					when "000100001111110" => rgb <= "000111";
					when "000100001111111" => rgb <= "000000";
					when "000100010000000" => rgb <= "101111";
					when "000100010000001" => rgb <= "000000";
					when "000100010000010" => rgb <= "000111";
					when "000100010000011" => rgb <= "000111";
					when "000100010000100" => rgb <= "000000";
					when "000100010000101" => rgb <= "000000";
					when "000100010000110" => rgb <= "000111";
					when "000100010000111" => rgb <= "000111";
					when "000100010001000" => rgb <= "000000";
					when "000100010001001" => rgb <= "101111";
					when "000100010001010" => rgb <= "000000";
					when "000100010001011" => rgb <= "000111";
					when "000100010001100" => rgb <= "000000";
					when "000100010001101" => rgb <= "000000";
					when "000100010001110" => rgb <= "000111";
					when "000100010001111" => rgb <= "000111";
					when "000100010010000" => rgb <= "000000";
					when "000100010010001" => rgb <= "101111";
					when "000100010010010" => rgb <= "000000";
					when "000100010010011" => rgb <= "000111";
					when "000100010010100" => rgb <= "000111";
					when "000100010010101" => rgb <= "000111";
					when "000100010010110" => rgb <= "000111";
					when "000100010010111" => rgb <= "000000";
					when "000100010011000" => rgb <= "101111";
					when "000100010011001" => rgb <= "000000";
					when "000100010011010" => rgb <= "000111";
					when "000100010011011" => rgb <= "000111";
					when "000100010011100" => rgb <= "000000";
					when "000100010011101" => rgb <= "101111";
					when "000100010011110" => rgb <= "101111";
					when "000100010011111" => rgb <= "101111";
					when "000100100000000" => rgb <= "101111";
					when "000100100000001" => rgb <= "101111";
					when "000100100000010" => rgb <= "101111";
					when "000100100000011" => rgb <= "101111";
					when "000100100000100" => rgb <= "101111";
					when "000100100000101" => rgb <= "101111";
					when "000100100000110" => rgb <= "000000";
					when "000100100000111" => rgb <= "000000";
					when "000100100001000" => rgb <= "000000";
					when "000100100001001" => rgb <= "110000";
					when "000100100001010" => rgb <= "110000";
					when "000100100001011" => rgb <= "000000";
					when "000100100001100" => rgb <= "000000";
					when "000100100001101" => rgb <= "000000";
					when "000100100001110" => rgb <= "101111";
					when "000100100001111" => rgb <= "000000";
					when "000100100010000" => rgb <= "110000";
					when "000100100010001" => rgb <= "110000";
					when "000100100010010" => rgb <= "000000";
					when "000100100010011" => rgb <= "110000";
					when "000100100010100" => rgb <= "110000";
					when "000100100010101" => rgb <= "000000";
					when "000100100010110" => rgb <= "101111";
					when "000100100010111" => rgb <= "000000";
					when "000100100011000" => rgb <= "110000";
					when "000100100011001" => rgb <= "110000";
					when "000100100011010" => rgb <= "000000";
					when "000100100011011" => rgb <= "110000";
					when "000100100011100" => rgb <= "110000";
					when "000100100011101" => rgb <= "000000";
					when "000100100011110" => rgb <= "101111";
					when "000100100011111" => rgb <= "000000";
					when "000100100100000" => rgb <= "110000";
					when "000100100100001" => rgb <= "110000";
					when "000100100100010" => rgb <= "110000";
					when "000100100100011" => rgb <= "110000";
					when "000100100100100" => rgb <= "110000";
					when "000100100100101" => rgb <= "110000";
					when "000100100100110" => rgb <= "000000";
					when "000100100100111" => rgb <= "101111";
					when "000100100101000" => rgb <= "000000";
					when "000100100101001" => rgb <= "000000";
					when "000100100101010" => rgb <= "101111";
					when "000100100101011" => rgb <= "101111";
					when "000100100101100" => rgb <= "101111";
					when "000100100101101" => rgb <= "101111";
					when "000100100101110" => rgb <= "101111";
					when "000100100101111" => rgb <= "101111";
					when "000100100110000" => rgb <= "101111";
					when "000100100110001" => rgb <= "101111";
					when "000100100110010" => rgb <= "101111";
					when "000100100110011" => rgb <= "101111";
					when "000100100110100" => rgb <= "101111";
					when "000100100110101" => rgb <= "101111";
					when "000100100110110" => rgb <= "101111";
					when "000100100110111" => rgb <= "101111";
					when "000100100111000" => rgb <= "101111";
					when "000100100111001" => rgb <= "101111";
					when "000100100111010" => rgb <= "101111";
					when "000100100111011" => rgb <= "101111";
					when "000100100111100" => rgb <= "101111";
					when "000100100111101" => rgb <= "101111";
					when "000100100111110" => rgb <= "101111";
					when "000100100111111" => rgb <= "101111";
					when "000100101000000" => rgb <= "101111";
					when "000100101000001" => rgb <= "101111";
					when "000100101000010" => rgb <= "101111";
					when "000100101000011" => rgb <= "101111";
					when "000100101000100" => rgb <= "101111";
					when "000100101000101" => rgb <= "101111";
					when "000100101000110" => rgb <= "101111";
					when "000100101000111" => rgb <= "101111";
					when "000100101001000" => rgb <= "101111";
					when "000100101001001" => rgb <= "101111";
					when "000100101001010" => rgb <= "101111";
					when "000100101001011" => rgb <= "101111";
					when "000100101001100" => rgb <= "101111";
					when "000100101001101" => rgb <= "101111";
					when "000100101001110" => rgb <= "101111";
					when "000100101001111" => rgb <= "101111";
					when "000100101010000" => rgb <= "101111";
					when "000100101010001" => rgb <= "101111";
					when "000100101010010" => rgb <= "101111";
					when "000100101010011" => rgb <= "101111";
					when "000100101010100" => rgb <= "101111";
					when "000100101010101" => rgb <= "101111";
					when "000100101010110" => rgb <= "101111";
					when "000100101010111" => rgb <= "101111";
					when "000100101011000" => rgb <= "101111";
					when "000100101011001" => rgb <= "101111";
					when "000100101011010" => rgb <= "101111";
					when "000100101011011" => rgb <= "101111";
					when "000100101011100" => rgb <= "101111";
					when "000100101011101" => rgb <= "101111";
					when "000100101011110" => rgb <= "101111";
					when "000100101011111" => rgb <= "101111";
					when "000100101100000" => rgb <= "101111";
					when "000100101100001" => rgb <= "101111";
					when "000100101100010" => rgb <= "101111";
					when "000100101100011" => rgb <= "101111";
					when "000100101100100" => rgb <= "101111";
					when "000100101100101" => rgb <= "101111";
					when "000100101100110" => rgb <= "101111";
					when "000100101100111" => rgb <= "101111";
					when "000100101101000" => rgb <= "101111";
					when "000100101101001" => rgb <= "101111";
					when "000100101101010" => rgb <= "101111";
					when "000100101101011" => rgb <= "101111";
					when "000100101101100" => rgb <= "101111";
					when "000100101101101" => rgb <= "101111";
					when "000100101101110" => rgb <= "101111";
					when "000100101101111" => rgb <= "101111";
					when "000100101110000" => rgb <= "101111";
					when "000100101110001" => rgb <= "101111";
					when "000100101110010" => rgb <= "101111";
					when "000100101110011" => rgb <= "101111";
					when "000100101110100" => rgb <= "101111";
					when "000100101110101" => rgb <= "101111";
					when "000100101110110" => rgb <= "000000";
					when "000100101110111" => rgb <= "000000";
					when "000100101111000" => rgb <= "101111";
					when "000100101111001" => rgb <= "000000";
					when "000100101111010" => rgb <= "000111";
					when "000100101111011" => rgb <= "000111";
					when "000100101111100" => rgb <= "000000";
					when "000100101111101" => rgb <= "000000";
					when "000100101111110" => rgb <= "000000";
					when "000100101111111" => rgb <= "000000";
					when "000100110000000" => rgb <= "101111";
					when "000100110000001" => rgb <= "000000";
					when "000100110000010" => rgb <= "000111";
					when "000100110000011" => rgb <= "000111";
					when "000100110000100" => rgb <= "000000";
					when "000100110000101" => rgb <= "000000";
					when "000100110000110" => rgb <= "000111";
					when "000100110000111" => rgb <= "000111";
					when "000100110001000" => rgb <= "000000";
					when "000100110001001" => rgb <= "101111";
					when "000100110001010" => rgb <= "000000";
					when "000100110001011" => rgb <= "000111";
					when "000100110001100" => rgb <= "000111";
					when "000100110001101" => rgb <= "000000";
					when "000100110001110" => rgb <= "000111";
					when "000100110001111" => rgb <= "000111";
					when "000100110010000" => rgb <= "000000";
					when "000100110010001" => rgb <= "101111";
					when "000100110010010" => rgb <= "000000";
					when "000100110010011" => rgb <= "000000";
					when "000100110010100" => rgb <= "000111";
					when "000100110010101" => rgb <= "000111";
					when "000100110010110" => rgb <= "000000";
					when "000100110010111" => rgb <= "000000";
					when "000100110011000" => rgb <= "101111";
					when "000100110011001" => rgb <= "000000";
					when "000100110011010" => rgb <= "000111";
					when "000100110011011" => rgb <= "000111";
					when "000100110011100" => rgb <= "000000";
					when "000100110011101" => rgb <= "101111";
					when "000100110011110" => rgb <= "101111";
					when "000100110011111" => rgb <= "101111";
					when "000101000000000" => rgb <= "101111";
					when "000101000000001" => rgb <= "101111";
					when "000101000000010" => rgb <= "101111";
					when "000101000000011" => rgb <= "101111";
					when "000101000000100" => rgb <= "101111";
					when "000101000000101" => rgb <= "101111";
					when "000101000000110" => rgb <= "101111";
					when "000101000000111" => rgb <= "101111";
					when "000101000001000" => rgb <= "000000";
					when "000101000001001" => rgb <= "100000";
					when "000101000001010" => rgb <= "100000";
					when "000101000001011" => rgb <= "000000";
					when "000101000001100" => rgb <= "000000";
					when "000101000001101" => rgb <= "101111";
					when "000101000001110" => rgb <= "101111";
					when "000101000001111" => rgb <= "000000";
					when "000101000010000" => rgb <= "100000";
					when "000101000010001" => rgb <= "100000";
					when "000101000010010" => rgb <= "000000";
					when "000101000010011" => rgb <= "100000";
					when "000101000010100" => rgb <= "100000";
					when "000101000010101" => rgb <= "000000";
					when "000101000010110" => rgb <= "101111";
					when "000101000010111" => rgb <= "000000";
					when "000101000011000" => rgb <= "100000";
					when "000101000011001" => rgb <= "100000";
					when "000101000011010" => rgb <= "100000";
					when "000101000011011" => rgb <= "100000";
					when "000101000011100" => rgb <= "100000";
					when "000101000011101" => rgb <= "000000";
					when "000101000011110" => rgb <= "101111";
					when "000101000011111" => rgb <= "000000";
					when "000101000100000" => rgb <= "000000";
					when "000101000100001" => rgb <= "100000";
					when "000101000100010" => rgb <= "100000";
					when "000101000100011" => rgb <= "100000";
					when "000101000100100" => rgb <= "100000";
					when "000101000100101" => rgb <= "000000";
					when "000101000100110" => rgb <= "000000";
					when "000101000100111" => rgb <= "101111";
					when "000101000101000" => rgb <= "000000";
					when "000101000101001" => rgb <= "000000";
					when "000101000101010" => rgb <= "101111";
					when "000101000101011" => rgb <= "101111";
					when "000101000101100" => rgb <= "101111";
					when "000101000101101" => rgb <= "101111";
					when "000101000101110" => rgb <= "101111";
					when "000101000101111" => rgb <= "101111";
					when "000101000110000" => rgb <= "101111";
					when "000101000110001" => rgb <= "101111";
					when "000101000110010" => rgb <= "101111";
					when "000101000110011" => rgb <= "101111";
					when "000101000110100" => rgb <= "101111";
					when "000101000110101" => rgb <= "101111";
					when "000101000110110" => rgb <= "101111";
					when "000101000110111" => rgb <= "101111";
					when "000101000111000" => rgb <= "101111";
					when "000101000111001" => rgb <= "101111";
					when "000101000111010" => rgb <= "101111";
					when "000101000111011" => rgb <= "101111";
					when "000101000111100" => rgb <= "101111";
					when "000101000111101" => rgb <= "101111";
					when "000101000111110" => rgb <= "101111";
					when "000101000111111" => rgb <= "101111";
					when "000101001000000" => rgb <= "101111";
					when "000101001000001" => rgb <= "101111";
					when "000101001000010" => rgb <= "101111";
					when "000101001000011" => rgb <= "101111";
					when "000101001000100" => rgb <= "101111";
					when "000101001000101" => rgb <= "101111";
					when "000101001000110" => rgb <= "101111";
					when "000101001000111" => rgb <= "101111";
					when "000101001001000" => rgb <= "101111";
					when "000101001001001" => rgb <= "101111";
					when "000101001001010" => rgb <= "101111";
					when "000101001001011" => rgb <= "101111";
					when "000101001001100" => rgb <= "101111";
					when "000101001001101" => rgb <= "101111";
					when "000101001001110" => rgb <= "101111";
					when "000101001001111" => rgb <= "101111";
					when "000101001010000" => rgb <= "101111";
					when "000101001010001" => rgb <= "101111";
					when "000101001010010" => rgb <= "101111";
					when "000101001010011" => rgb <= "101111";
					when "000101001010100" => rgb <= "101111";
					when "000101001010101" => rgb <= "101111";
					when "000101001010110" => rgb <= "101111";
					when "000101001010111" => rgb <= "101111";
					when "000101001011000" => rgb <= "101111";
					when "000101001011001" => rgb <= "101111";
					when "000101001011010" => rgb <= "101111";
					when "000101001011011" => rgb <= "101111";
					when "000101001011100" => rgb <= "101111";
					when "000101001011101" => rgb <= "101111";
					when "000101001011110" => rgb <= "101111";
					when "000101001011111" => rgb <= "101111";
					when "000101001100000" => rgb <= "101111";
					when "000101001100001" => rgb <= "101111";
					when "000101001100010" => rgb <= "101111";
					when "000101001100011" => rgb <= "101111";
					when "000101001100100" => rgb <= "101111";
					when "000101001100101" => rgb <= "101111";
					when "000101001100110" => rgb <= "101111";
					when "000101001100111" => rgb <= "101111";
					when "000101001101000" => rgb <= "101111";
					when "000101001101001" => rgb <= "101111";
					when "000101001101010" => rgb <= "101111";
					when "000101001101011" => rgb <= "101111";
					when "000101001101100" => rgb <= "101111";
					when "000101001101101" => rgb <= "101111";
					when "000101001101110" => rgb <= "101111";
					when "000101001101111" => rgb <= "101111";
					when "000101001110000" => rgb <= "101111";
					when "000101001110001" => rgb <= "101111";
					when "000101001110010" => rgb <= "101111";
					when "000101001110011" => rgb <= "101111";
					when "000101001110100" => rgb <= "101111";
					when "000101001110101" => rgb <= "101111";
					when "000101001110110" => rgb <= "000000";
					when "000101001110111" => rgb <= "000000";
					when "000101001111000" => rgb <= "101111";
					when "000101001111001" => rgb <= "000000";
					when "000101001111010" => rgb <= "000000";
					when "000101001111011" => rgb <= "000110";
					when "000101001111100" => rgb <= "000110";
					when "000101001111101" => rgb <= "000110";
					when "000101001111110" => rgb <= "000110";
					when "000101001111111" => rgb <= "000000";
					when "000101010000000" => rgb <= "101111";
					when "000101010000001" => rgb <= "000000";
					when "000101010000010" => rgb <= "000110";
					when "000101010000011" => rgb <= "000110";
					when "000101010000100" => rgb <= "000000";
					when "000101010000101" => rgb <= "000000";
					when "000101010000110" => rgb <= "000110";
					when "000101010000111" => rgb <= "000110";
					when "000101010001000" => rgb <= "000000";
					when "000101010001001" => rgb <= "101111";
					when "000101010001010" => rgb <= "000000";
					when "000101010001011" => rgb <= "000110";
					when "000101010001100" => rgb <= "000110";
					when "000101010001101" => rgb <= "000110";
					when "000101010001110" => rgb <= "000110";
					when "000101010001111" => rgb <= "000110";
					when "000101010010000" => rgb <= "000000";
					when "000101010010001" => rgb <= "101111";
					when "000101010010010" => rgb <= "101111";
					when "000101010010011" => rgb <= "000000";
					when "000101010010100" => rgb <= "000110";
					when "000101010010101" => rgb <= "000110";
					when "000101010010110" => rgb <= "000000";
					when "000101010010111" => rgb <= "101111";
					when "000101010011000" => rgb <= "101111";
					when "000101010011001" => rgb <= "000000";
					when "000101010011010" => rgb <= "000110";
					when "000101010011011" => rgb <= "000110";
					when "000101010011100" => rgb <= "000000";
					when "000101010011101" => rgb <= "101111";
					when "000101010011110" => rgb <= "101111";
					when "000101010011111" => rgb <= "101111";
					when "000101100000000" => rgb <= "101111";
					when "000101100000001" => rgb <= "101111";
					when "000101100000010" => rgb <= "101111";
					when "000101100000011" => rgb <= "101111";
					when "000101100000100" => rgb <= "101111";
					when "000101100000101" => rgb <= "101111";
					when "000101100000110" => rgb <= "000000";
					when "000101100000111" => rgb <= "101111";
					when "000101100001000" => rgb <= "000000";
					when "000101100001001" => rgb <= "100000";
					when "000101100001010" => rgb <= "100000";
					when "000101100001011" => rgb <= "000000";
					when "000101100001100" => rgb <= "101111";
					when "000101100001101" => rgb <= "001000";
					when "000101100001110" => rgb <= "101111";
					when "000101100001111" => rgb <= "000000";
					when "000101100010000" => rgb <= "100000";
					when "000101100010001" => rgb <= "100000";
					when "000101100010010" => rgb <= "000000";
					when "000101100010011" => rgb <= "100000";
					when "000101100010100" => rgb <= "100000";
					when "000101100010101" => rgb <= "000000";
					when "000101100010110" => rgb <= "101111";
					when "000101100010111" => rgb <= "000000";
					when "000101100011000" => rgb <= "100000";
					when "000101100011001" => rgb <= "100000";
					when "000101100011010" => rgb <= "000000";
					when "000101100011011" => rgb <= "100000";
					when "000101100011100" => rgb <= "100000";
					when "000101100011101" => rgb <= "000000";
					when "000101100011110" => rgb <= "101111";
					when "000101100011111" => rgb <= "101111";
					when "000101100100000" => rgb <= "000000";
					when "000101100100001" => rgb <= "000000";
					when "000101100100010" => rgb <= "100000";
					when "000101100100011" => rgb <= "100000";
					when "000101100100100" => rgb <= "000000";
					when "000101100100101" => rgb <= "000000";
					when "000101100100110" => rgb <= "101111";
					when "000101100100111" => rgb <= "101111";
					when "000101100101000" => rgb <= "000000";
					when "000101100101001" => rgb <= "000000";
					when "000101100101010" => rgb <= "101111";
					when "000101100101011" => rgb <= "101111";
					when "000101100101100" => rgb <= "101111";
					when "000101100101101" => rgb <= "101111";
					when "000101100101110" => rgb <= "101111";
					when "000101100101111" => rgb <= "101111";
					when "000101100110000" => rgb <= "101111";
					when "000101100110001" => rgb <= "101111";
					when "000101100110010" => rgb <= "101111";
					when "000101100110011" => rgb <= "101111";
					when "000101100110100" => rgb <= "101111";
					when "000101100110101" => rgb <= "101111";
					when "000101100110110" => rgb <= "101111";
					when "000101100110111" => rgb <= "101111";
					when "000101100111000" => rgb <= "101111";
					when "000101100111001" => rgb <= "101111";
					when "000101100111010" => rgb <= "101111";
					when "000101100111011" => rgb <= "101111";
					when "000101100111100" => rgb <= "101111";
					when "000101100111101" => rgb <= "101111";
					when "000101100111110" => rgb <= "101111";
					when "000101100111111" => rgb <= "101111";
					when "000101101000000" => rgb <= "101111";
					when "000101101000001" => rgb <= "101111";
					when "000101101000010" => rgb <= "101111";
					when "000101101000011" => rgb <= "101111";
					when "000101101000100" => rgb <= "101111";
					when "000101101000101" => rgb <= "101111";
					when "000101101000110" => rgb <= "101111";
					when "000101101000111" => rgb <= "101111";
					when "000101101001000" => rgb <= "101111";
					when "000101101001001" => rgb <= "101111";
					when "000101101001010" => rgb <= "101111";
					when "000101101001011" => rgb <= "101111";
					when "000101101001100" => rgb <= "101111";
					when "000101101001101" => rgb <= "101111";
					when "000101101001110" => rgb <= "101111";
					when "000101101001111" => rgb <= "101111";
					when "000101101010000" => rgb <= "101111";
					when "000101101010001" => rgb <= "101111";
					when "000101101010010" => rgb <= "101111";
					when "000101101010011" => rgb <= "101111";
					when "000101101010100" => rgb <= "101111";
					when "000101101010101" => rgb <= "101111";
					when "000101101010110" => rgb <= "101111";
					when "000101101010111" => rgb <= "101111";
					when "000101101011000" => rgb <= "101111";
					when "000101101011001" => rgb <= "101111";
					when "000101101011010" => rgb <= "101111";
					when "000101101011011" => rgb <= "101111";
					when "000101101011100" => rgb <= "101111";
					when "000101101011101" => rgb <= "101111";
					when "000101101011110" => rgb <= "101111";
					when "000101101011111" => rgb <= "101111";
					when "000101101100000" => rgb <= "101111";
					when "000101101100001" => rgb <= "101111";
					when "000101101100010" => rgb <= "101111";
					when "000101101100011" => rgb <= "101111";
					when "000101101100100" => rgb <= "101111";
					when "000101101100101" => rgb <= "101111";
					when "000101101100110" => rgb <= "101111";
					when "000101101100111" => rgb <= "101111";
					when "000101101101000" => rgb <= "101111";
					when "000101101101001" => rgb <= "101111";
					when "000101101101010" => rgb <= "101111";
					when "000101101101011" => rgb <= "101111";
					when "000101101101100" => rgb <= "101111";
					when "000101101101101" => rgb <= "101111";
					when "000101101101110" => rgb <= "101111";
					when "000101101101111" => rgb <= "101111";
					when "000101101110000" => rgb <= "101111";
					when "000101101110001" => rgb <= "101111";
					when "000101101110010" => rgb <= "101111";
					when "000101101110011" => rgb <= "101111";
					when "000101101110100" => rgb <= "101111";
					when "000101101110101" => rgb <= "101111";
					when "000101101110110" => rgb <= "000000";
					when "000101101110111" => rgb <= "000000";
					when "000101101111000" => rgb <= "101111";
					when "000101101111001" => rgb <= "000000";
					when "000101101111010" => rgb <= "000000";
					when "000101101111011" => rgb <= "000000";
					when "000101101111100" => rgb <= "000000";
					when "000101101111101" => rgb <= "000110";
					when "000101101111110" => rgb <= "000110";
					when "000101101111111" => rgb <= "000000";
					when "000101110000000" => rgb <= "101111";
					when "000101110000001" => rgb <= "000000";
					when "000101110000010" => rgb <= "000110";
					when "000101110000011" => rgb <= "000110";
					when "000101110000100" => rgb <= "000000";
					when "000101110000101" => rgb <= "000000";
					when "000101110000110" => rgb <= "000110";
					when "000101110000111" => rgb <= "000110";
					when "000101110001000" => rgb <= "000000";
					when "000101110001001" => rgb <= "101111";
					when "000101110001010" => rgb <= "000000";
					when "000101110001011" => rgb <= "000110";
					when "000101110001100" => rgb <= "000110";
					when "000101110001101" => rgb <= "000000";
					when "000101110001110" => rgb <= "000110";
					when "000101110001111" => rgb <= "000110";
					when "000101110010000" => rgb <= "000000";
					when "000101110010001" => rgb <= "101111";
					when "000101110010010" => rgb <= "101111";
					when "000101110010011" => rgb <= "000000";
					when "000101110010100" => rgb <= "000110";
					when "000101110010101" => rgb <= "000110";
					when "000101110010110" => rgb <= "000000";
					when "000101110010111" => rgb <= "101111";
					when "000101110011000" => rgb <= "101111";
					when "000101110011001" => rgb <= "000000";
					when "000101110011010" => rgb <= "000110";
					when "000101110011011" => rgb <= "000110";
					when "000101110011100" => rgb <= "000000";
					when "000101110011101" => rgb <= "000000";
					when "000101110011110" => rgb <= "101111";
					when "000101110011111" => rgb <= "101111";
					when "000110000000000" => rgb <= "101111";
					when "000110000000001" => rgb <= "101111";
					when "000110000000010" => rgb <= "101111";
					when "000110000000011" => rgb <= "101111";
					when "000110000000100" => rgb <= "101111";
					when "000110000000101" => rgb <= "101111";
					when "000110000000110" => rgb <= "000000";
					when "000110000000111" => rgb <= "101111";
					when "000110000001000" => rgb <= "000000";
					when "000110000001001" => rgb <= "010000";
					when "000110000001010" => rgb <= "010000";
					when "000110000001011" => rgb <= "000000";
					when "000110000001100" => rgb <= "101111";
					when "000110000001101" => rgb <= "001000";
					when "000110000001110" => rgb <= "101111";
					when "000110000001111" => rgb <= "000000";
					when "000110000010000" => rgb <= "000000";
					when "000110000010001" => rgb <= "010000";
					when "000110000010010" => rgb <= "010000";
					when "000110000010011" => rgb <= "010000";
					when "000110000010100" => rgb <= "000000";
					when "000110000010101" => rgb <= "000000";
					when "000110000010110" => rgb <= "101111";
					when "000110000010111" => rgb <= "000000";
					when "000110000011000" => rgb <= "010000";
					when "000110000011001" => rgb <= "010000";
					when "000110000011010" => rgb <= "000000";
					when "000110000011011" => rgb <= "010000";
					when "000110000011100" => rgb <= "010000";
					when "000110000011101" => rgb <= "000000";
					when "000110000011110" => rgb <= "101111";
					when "000110000011111" => rgb <= "101111";
					when "000110000100000" => rgb <= "101111";
					when "000110000100001" => rgb <= "000000";
					when "000110000100010" => rgb <= "010000";
					when "000110000100011" => rgb <= "010000";
					when "000110000100100" => rgb <= "000000";
					when "000110000100101" => rgb <= "101111";
					when "000110000100110" => rgb <= "101111";
					when "000110000100111" => rgb <= "001000";
					when "000110000101000" => rgb <= "000000";
					when "000110000101001" => rgb <= "000000";
					when "000110000101010" => rgb <= "101111";
					when "000110000101011" => rgb <= "101111";
					when "000110000101100" => rgb <= "101111";
					when "000110000101101" => rgb <= "101111";
					when "000110000101110" => rgb <= "101111";
					when "000110000101111" => rgb <= "101111";
					when "000110000110000" => rgb <= "101111";
					when "000110000110001" => rgb <= "101111";
					when "000110000110010" => rgb <= "101111";
					when "000110000110011" => rgb <= "101111";
					when "000110000110100" => rgb <= "101111";
					when "000110000110101" => rgb <= "101111";
					when "000110000110110" => rgb <= "101111";
					when "000110000110111" => rgb <= "101111";
					when "000110000111000" => rgb <= "101111";
					when "000110000111001" => rgb <= "101111";
					when "000110000111010" => rgb <= "101111";
					when "000110000111011" => rgb <= "101111";
					when "000110000111100" => rgb <= "101111";
					when "000110000111101" => rgb <= "101111";
					when "000110000111110" => rgb <= "101111";
					when "000110000111111" => rgb <= "101111";
					when "000110001000000" => rgb <= "101111";
					when "000110001000001" => rgb <= "101111";
					when "000110001000010" => rgb <= "101111";
					when "000110001000011" => rgb <= "101111";
					when "000110001000100" => rgb <= "101111";
					when "000110001000101" => rgb <= "101111";
					when "000110001000110" => rgb <= "101111";
					when "000110001000111" => rgb <= "101111";
					when "000110001001000" => rgb <= "101111";
					when "000110001001001" => rgb <= "101111";
					when "000110001001010" => rgb <= "101111";
					when "000110001001011" => rgb <= "101111";
					when "000110001001100" => rgb <= "101111";
					when "000110001001101" => rgb <= "101111";
					when "000110001001110" => rgb <= "101111";
					when "000110001001111" => rgb <= "101111";
					when "000110001010000" => rgb <= "101111";
					when "000110001010001" => rgb <= "101111";
					when "000110001010010" => rgb <= "101111";
					when "000110001010011" => rgb <= "101111";
					when "000110001010100" => rgb <= "101111";
					when "000110001010101" => rgb <= "101111";
					when "000110001010110" => rgb <= "101111";
					when "000110001010111" => rgb <= "101111";
					when "000110001011000" => rgb <= "101111";
					when "000110001011001" => rgb <= "101111";
					when "000110001011010" => rgb <= "101111";
					when "000110001011011" => rgb <= "101111";
					when "000110001011100" => rgb <= "101111";
					when "000110001011101" => rgb <= "101111";
					when "000110001011110" => rgb <= "101111";
					when "000110001011111" => rgb <= "101111";
					when "000110001100000" => rgb <= "101111";
					when "000110001100001" => rgb <= "101111";
					when "000110001100010" => rgb <= "101111";
					when "000110001100011" => rgb <= "101111";
					when "000110001100100" => rgb <= "101111";
					when "000110001100101" => rgb <= "101111";
					when "000110001100110" => rgb <= "101111";
					when "000110001100111" => rgb <= "101111";
					when "000110001101000" => rgb <= "101111";
					when "000110001101001" => rgb <= "101111";
					when "000110001101010" => rgb <= "101111";
					when "000110001101011" => rgb <= "101111";
					when "000110001101100" => rgb <= "101111";
					when "000110001101101" => rgb <= "101111";
					when "000110001101110" => rgb <= "101111";
					when "000110001101111" => rgb <= "101111";
					when "000110001110000" => rgb <= "101111";
					when "000110001110001" => rgb <= "101111";
					when "000110001110010" => rgb <= "101111";
					when "000110001110011" => rgb <= "101111";
					when "000110001110100" => rgb <= "101111";
					when "000110001110101" => rgb <= "101111";
					when "000110001110110" => rgb <= "000000";
					when "000110001110111" => rgb <= "000000";
					when "000110001111000" => rgb <= "101111";
					when "000110001111001" => rgb <= "000000";
					when "000110001111010" => rgb <= "000011";
					when "000110001111011" => rgb <= "000011";
					when "000110001111100" => rgb <= "000011";
					when "000110001111101" => rgb <= "000011";
					when "000110001111110" => rgb <= "000011";
					when "000110001111111" => rgb <= "000000";
					when "000110010000000" => rgb <= "101111";
					when "000110010000001" => rgb <= "000000";
					when "000110010000010" => rgb <= "000000";
					when "000110010000011" => rgb <= "000011";
					when "000110010000100" => rgb <= "000011";
					when "000110010000101" => rgb <= "000011";
					when "000110010000110" => rgb <= "000011";
					when "000110010000111" => rgb <= "000000";
					when "000110010001000" => rgb <= "000000";
					when "000110010001001" => rgb <= "101111";
					when "000110010001010" => rgb <= "000000";
					when "000110010001011" => rgb <= "000011";
					when "000110010001100" => rgb <= "000011";
					when "000110010001101" => rgb <= "000000";
					when "000110010001110" => rgb <= "000011";
					when "000110010001111" => rgb <= "000011";
					when "000110010010000" => rgb <= "000000";
					when "000110010010001" => rgb <= "101111";
					when "000110010010010" => rgb <= "000000";
					when "000110010010011" => rgb <= "000011";
					when "000110010010100" => rgb <= "000011";
					when "000110010010101" => rgb <= "000011";
					when "000110010010110" => rgb <= "000011";
					when "000110010010111" => rgb <= "000000";
					when "000110010011000" => rgb <= "101111";
					when "000110010011001" => rgb <= "000000";
					when "000110010011010" => rgb <= "000011";
					when "000110010011011" => rgb <= "000011";
					when "000110010011100" => rgb <= "000011";
					when "000110010011101" => rgb <= "000011";
					when "000110010011110" => rgb <= "000000";
					when "000110010011111" => rgb <= "101111";
					when "000110100000000" => rgb <= "101111";
					when "000110100000001" => rgb <= "101111";
					when "000110100000010" => rgb <= "101111";
					when "000110100000011" => rgb <= "101111";
					when "000110100000100" => rgb <= "101111";
					when "000110100000101" => rgb <= "101111";
					when "000110100000110" => rgb <= "000000";
					when "000110100000111" => rgb <= "101111";
					when "000110100001000" => rgb <= "000000";
					when "000110100001001" => rgb <= "000000";
					when "000110100001010" => rgb <= "000000";
					when "000110100001011" => rgb <= "000000";
					when "000110100001100" => rgb <= "101111";
					when "000110100001101" => rgb <= "001000";
					when "000110100001110" => rgb <= "101111";
					when "000110100001111" => rgb <= "101111";
					when "000110100010000" => rgb <= "000000";
					when "000110100010001" => rgb <= "000000";
					when "000110100010010" => rgb <= "000000";
					when "000110100010011" => rgb <= "000000";
					when "000110100010100" => rgb <= "000000";
					when "000110100010101" => rgb <= "101111";
					when "000110100010110" => rgb <= "101111";
					when "000110100010111" => rgb <= "000000";
					when "000110100011000" => rgb <= "000000";
					when "000110100011001" => rgb <= "000000";
					when "000110100011010" => rgb <= "000000";
					when "000110100011011" => rgb <= "000000";
					when "000110100011100" => rgb <= "000000";
					when "000110100011101" => rgb <= "000000";
					when "000110100011110" => rgb <= "101111";
					when "000110100011111" => rgb <= "001000";
					when "000110100100000" => rgb <= "101111";
					when "000110100100001" => rgb <= "000000";
					when "000110100100010" => rgb <= "000000";
					when "000110100100011" => rgb <= "000000";
					when "000110100100100" => rgb <= "000000";
					when "000110100100101" => rgb <= "101111";
					when "000110100100110" => rgb <= "001000";
					when "000110100100111" => rgb <= "001000";
					when "000110100101000" => rgb <= "000000";
					when "000110100101001" => rgb <= "000000";
					when "000110100101010" => rgb <= "101111";
					when "000110100101011" => rgb <= "101111";
					when "000110100101100" => rgb <= "101111";
					when "000110100101101" => rgb <= "101111";
					when "000110100101110" => rgb <= "101111";
					when "000110100101111" => rgb <= "101111";
					when "000110100110000" => rgb <= "101111";
					when "000110100110001" => rgb <= "101111";
					when "000110100110010" => rgb <= "101111";
					when "000110100110011" => rgb <= "101111";
					when "000110100110100" => rgb <= "101111";
					when "000110100110101" => rgb <= "101111";
					when "000110100110110" => rgb <= "101111";
					when "000110100110111" => rgb <= "101111";
					when "000110100111000" => rgb <= "101111";
					when "000110100111001" => rgb <= "101111";
					when "000110100111010" => rgb <= "101111";
					when "000110100111011" => rgb <= "101111";
					when "000110100111100" => rgb <= "101111";
					when "000110100111101" => rgb <= "101111";
					when "000110100111110" => rgb <= "101111";
					when "000110100111111" => rgb <= "101111";
					when "000110101000000" => rgb <= "101111";
					when "000110101000001" => rgb <= "101111";
					when "000110101000010" => rgb <= "101111";
					when "000110101000011" => rgb <= "101111";
					when "000110101000100" => rgb <= "101111";
					when "000110101000101" => rgb <= "101111";
					when "000110101000110" => rgb <= "101111";
					when "000110101000111" => rgb <= "101111";
					when "000110101001000" => rgb <= "101111";
					when "000110101001001" => rgb <= "101111";
					when "000110101001010" => rgb <= "101111";
					when "000110101001011" => rgb <= "101111";
					when "000110101001100" => rgb <= "101111";
					when "000110101001101" => rgb <= "101111";
					when "000110101001110" => rgb <= "101111";
					when "000110101001111" => rgb <= "101111";
					when "000110101010000" => rgb <= "101111";
					when "000110101010001" => rgb <= "101111";
					when "000110101010010" => rgb <= "101111";
					when "000110101010011" => rgb <= "101111";
					when "000110101010100" => rgb <= "101111";
					when "000110101010101" => rgb <= "101111";
					when "000110101010110" => rgb <= "101111";
					when "000110101010111" => rgb <= "101111";
					when "000110101011000" => rgb <= "101111";
					when "000110101011001" => rgb <= "101111";
					when "000110101011010" => rgb <= "101111";
					when "000110101011011" => rgb <= "101111";
					when "000110101011100" => rgb <= "101111";
					when "000110101011101" => rgb <= "101111";
					when "000110101011110" => rgb <= "101111";
					when "000110101011111" => rgb <= "101111";
					when "000110101100000" => rgb <= "101111";
					when "000110101100001" => rgb <= "101111";
					when "000110101100010" => rgb <= "101111";
					when "000110101100011" => rgb <= "101111";
					when "000110101100100" => rgb <= "101111";
					when "000110101100101" => rgb <= "101111";
					when "000110101100110" => rgb <= "101111";
					when "000110101100111" => rgb <= "101111";
					when "000110101101000" => rgb <= "101111";
					when "000110101101001" => rgb <= "101111";
					when "000110101101010" => rgb <= "101111";
					when "000110101101011" => rgb <= "101111";
					when "000110101101100" => rgb <= "101111";
					when "000110101101101" => rgb <= "101111";
					when "000110101101110" => rgb <= "101111";
					when "000110101101111" => rgb <= "101111";
					when "000110101110000" => rgb <= "101111";
					when "000110101110001" => rgb <= "101111";
					when "000110101110010" => rgb <= "101111";
					when "000110101110011" => rgb <= "101111";
					when "000110101110100" => rgb <= "101111";
					when "000110101110101" => rgb <= "101111";
					when "000110101110110" => rgb <= "000000";
					when "000110101110111" => rgb <= "000000";
					when "000110101111000" => rgb <= "101111";
					when "000110101111001" => rgb <= "000000";
					when "000110101111010" => rgb <= "000000";
					when "000110101111011" => rgb <= "000000";
					when "000110101111100" => rgb <= "000000";
					when "000110101111101" => rgb <= "000000";
					when "000110101111110" => rgb <= "000000";
					when "000110101111111" => rgb <= "101111";
					when "000110110000000" => rgb <= "101111";
					when "000110110000001" => rgb <= "101111";
					when "000110110000010" => rgb <= "000000";
					when "000110110000011" => rgb <= "000000";
					when "000110110000100" => rgb <= "000000";
					when "000110110000101" => rgb <= "000000";
					when "000110110000110" => rgb <= "000000";
					when "000110110000111" => rgb <= "000000";
					when "000110110001000" => rgb <= "101111";
					when "000110110001001" => rgb <= "101111";
					when "000110110001010" => rgb <= "000000";
					when "000110110001011" => rgb <= "000000";
					when "000110110001100" => rgb <= "000000";
					when "000110110001101" => rgb <= "000000";
					when "000110110001110" => rgb <= "000000";
					when "000110110001111" => rgb <= "000000";
					when "000110110010000" => rgb <= "000000";
					when "000110110010001" => rgb <= "101111";
					when "000110110010010" => rgb <= "000000";
					when "000110110010011" => rgb <= "000000";
					when "000110110010100" => rgb <= "000000";
					when "000110110010101" => rgb <= "000000";
					when "000110110010110" => rgb <= "000000";
					when "000110110010111" => rgb <= "000000";
					when "000110110011000" => rgb <= "101111";
					when "000110110011001" => rgb <= "000000";
					when "000110110011010" => rgb <= "000000";
					when "000110110011011" => rgb <= "000000";
					when "000110110011100" => rgb <= "000000";
					when "000110110011101" => rgb <= "000000";
					when "000110110011110" => rgb <= "000000";
					when "000110110011111" => rgb <= "101111";
					when "000111000000000" => rgb <= "101111";
					when "000111000000001" => rgb <= "101111";
					when "000111000000010" => rgb <= "101111";
					when "000111000000011" => rgb <= "101111";
					when "000111000000100" => rgb <= "000000";
					when "000111000000101" => rgb <= "000000";
					when "000111000000110" => rgb <= "001000";
					when "000111000000111" => rgb <= "101111";
					when "000111000001000" => rgb <= "101111";
					when "000111000001001" => rgb <= "000000";
					when "000111000001010" => rgb <= "000000";
					when "000111000001011" => rgb <= "101111";
					when "000111000001100" => rgb <= "101111";
					when "000111000001101" => rgb <= "001000";
					when "000111000001110" => rgb <= "001000";
					when "000111000001111" => rgb <= "101111";
					when "000111000010000" => rgb <= "101111";
					when "000111000010001" => rgb <= "000000";
					when "000111000010010" => rgb <= "000000";
					when "000111000010011" => rgb <= "000000";
					when "000111000010100" => rgb <= "101111";
					when "000111000010101" => rgb <= "101111";
					when "000111000010110" => rgb <= "001000";
					when "000111000010111" => rgb <= "101111";
					when "000111000011000" => rgb <= "000000";
					when "000111000011001" => rgb <= "000000";
					when "000111000011010" => rgb <= "101111";
					when "000111000011011" => rgb <= "000000";
					when "000111000011100" => rgb <= "000000";
					when "000111000011101" => rgb <= "101111";
					when "000111000011110" => rgb <= "101111";
					when "000111000011111" => rgb <= "001000";
					when "000111000100000" => rgb <= "101111";
					when "000111000100001" => rgb <= "101111";
					when "000111000100010" => rgb <= "000000";
					when "000111000100011" => rgb <= "000000";
					when "000111000100100" => rgb <= "101111";
					when "000111000100101" => rgb <= "101111";
					when "000111000100110" => rgb <= "001000";
					when "000111000100111" => rgb <= "001000";
					when "000111000101000" => rgb <= "000000";
					when "000111000101001" => rgb <= "000000";
					when "000111000101010" => rgb <= "000000";
					when "000111000101011" => rgb <= "000000";
					when "000111000101100" => rgb <= "000000";
					when "000111000101101" => rgb <= "000000";
					when "000111000101110" => rgb <= "000000";
					when "000111000101111" => rgb <= "000000";
					when "000111000110000" => rgb <= "000000";
					when "000111000110001" => rgb <= "000000";
					when "000111000110010" => rgb <= "000000";
					when "000111000110011" => rgb <= "000000";
					when "000111000110100" => rgb <= "000000";
					when "000111000110101" => rgb <= "000000";
					when "000111000110110" => rgb <= "000000";
					when "000111000110111" => rgb <= "000000";
					when "000111000111000" => rgb <= "000000";
					when "000111000111001" => rgb <= "000000";
					when "000111000111010" => rgb <= "000000";
					when "000111000111011" => rgb <= "000000";
					when "000111000111100" => rgb <= "000000";
					when "000111000111101" => rgb <= "000000";
					when "000111000111110" => rgb <= "000000";
					when "000111000111111" => rgb <= "000000";
					when "000111001000000" => rgb <= "000000";
					when "000111001000001" => rgb <= "000000";
					when "000111001000010" => rgb <= "000000";
					when "000111001000011" => rgb <= "000000";
					when "000111001000100" => rgb <= "000000";
					when "000111001000101" => rgb <= "000000";
					when "000111001000110" => rgb <= "000000";
					when "000111001000111" => rgb <= "000000";
					when "000111001001000" => rgb <= "000000";
					when "000111001001001" => rgb <= "000000";
					when "000111001001010" => rgb <= "000000";
					when "000111001001011" => rgb <= "000000";
					when "000111001001100" => rgb <= "000000";
					when "000111001001101" => rgb <= "000000";
					when "000111001001110" => rgb <= "000000";
					when "000111001001111" => rgb <= "000000";
					when "000111001010000" => rgb <= "000000";
					when "000111001010001" => rgb <= "000000";
					when "000111001010010" => rgb <= "000000";
					when "000111001010011" => rgb <= "000000";
					when "000111001010100" => rgb <= "000000";
					when "000111001010101" => rgb <= "000000";
					when "000111001010110" => rgb <= "000000";
					when "000111001010111" => rgb <= "000000";
					when "000111001011000" => rgb <= "000000";
					when "000111001011001" => rgb <= "000000";
					when "000111001011010" => rgb <= "000000";
					when "000111001011011" => rgb <= "000000";
					when "000111001011100" => rgb <= "000000";
					when "000111001011101" => rgb <= "000000";
					when "000111001011110" => rgb <= "000000";
					when "000111001011111" => rgb <= "000000";
					when "000111001100000" => rgb <= "000000";
					when "000111001100001" => rgb <= "000000";
					when "000111001100010" => rgb <= "000000";
					when "000111001100011" => rgb <= "000000";
					when "000111001100100" => rgb <= "000000";
					when "000111001100101" => rgb <= "000000";
					when "000111001100110" => rgb <= "000000";
					when "000111001100111" => rgb <= "000000";
					when "000111001101000" => rgb <= "000000";
					when "000111001101001" => rgb <= "000000";
					when "000111001101010" => rgb <= "000000";
					when "000111001101011" => rgb <= "000000";
					when "000111001101100" => rgb <= "000000";
					when "000111001101101" => rgb <= "000000";
					when "000111001101110" => rgb <= "000000";
					when "000111001101111" => rgb <= "000000";
					when "000111001110000" => rgb <= "000000";
					when "000111001110001" => rgb <= "000000";
					when "000111001110010" => rgb <= "000000";
					when "000111001110011" => rgb <= "000000";
					when "000111001110100" => rgb <= "000000";
					when "000111001110101" => rgb <= "000000";
					when "000111001110110" => rgb <= "000000";
					when "000111001110111" => rgb <= "000000";
					when "000111001111000" => rgb <= "101111";
					when "000111001111001" => rgb <= "101111";
					when "000111001111010" => rgb <= "000000";
					when "000111001111011" => rgb <= "000000";
					when "000111001111100" => rgb <= "000000";
					when "000111001111101" => rgb <= "000000";
					when "000111001111110" => rgb <= "101111";
					when "000111001111111" => rgb <= "101111";
					when "000111010000000" => rgb <= "101111";
					when "000111010000001" => rgb <= "101111";
					when "000111010000010" => rgb <= "101111";
					when "000111010000011" => rgb <= "000000";
					when "000111010000100" => rgb <= "000000";
					when "000111010000101" => rgb <= "000000";
					when "000111010000110" => rgb <= "000000";
					when "000111010000111" => rgb <= "101111";
					when "000111010001000" => rgb <= "101111";
					when "000111010001001" => rgb <= "101111";
					when "000111010001010" => rgb <= "101111";
					when "000111010001011" => rgb <= "000000";
					when "000111010001100" => rgb <= "000000";
					when "000111010001101" => rgb <= "101111";
					when "000111010001110" => rgb <= "000000";
					when "000111010001111" => rgb <= "000000";
					when "000111010010000" => rgb <= "101111";
					when "000111010010001" => rgb <= "101111";
					when "000111010010010" => rgb <= "101111";
					when "000111010010011" => rgb <= "000000";
					when "000111010010100" => rgb <= "000000";
					when "000111010010101" => rgb <= "000000";
					when "000111010010110" => rgb <= "000000";
					when "000111010010111" => rgb <= "101111";
					when "000111010011000" => rgb <= "101111";
					when "000111010011001" => rgb <= "101111";
					when "000111010011010" => rgb <= "000000";
					when "000111010011011" => rgb <= "000000";
					when "000111010011100" => rgb <= "000000";
					when "000111010011101" => rgb <= "000000";
					when "000111010011110" => rgb <= "101111";
					when "000111010011111" => rgb <= "101111";
					when "000111100000000" => rgb <= "101111";
					when "000111100000001" => rgb <= "101111";
					when "000111100000010" => rgb <= "101111";
					when "000111100000011" => rgb <= "101111";
					when "000111100000100" => rgb <= "000000";
					when "000111100000101" => rgb <= "000000";
					when "000111100000110" => rgb <= "001000";
					when "000111100000111" => rgb <= "001000";
					when "000111100001000" => rgb <= "101111";
					when "000111100001001" => rgb <= "101111";
					when "000111100001010" => rgb <= "101111";
					when "000111100001011" => rgb <= "101111";
					when "000111100001100" => rgb <= "001000";
					when "000111100001101" => rgb <= "001000";
					when "000111100001110" => rgb <= "001000";
					when "000111100001111" => rgb <= "001000";
					when "000111100010000" => rgb <= "101111";
					when "000111100010001" => rgb <= "101111";
					when "000111100010010" => rgb <= "101111";
					when "000111100010011" => rgb <= "101111";
					when "000111100010100" => rgb <= "101111";
					when "000111100010101" => rgb <= "001000";
					when "000111100010110" => rgb <= "001000";
					when "000111100010111" => rgb <= "101111";
					when "000111100011000" => rgb <= "101111";
					when "000111100011001" => rgb <= "101111";
					when "000111100011010" => rgb <= "101111";
					when "000111100011011" => rgb <= "101111";
					when "000111100011100" => rgb <= "101111";
					when "000111100011101" => rgb <= "101111";
					when "000111100011110" => rgb <= "001000";
					when "000111100011111" => rgb <= "001000";
					when "000111100100000" => rgb <= "001000";
					when "000111100100001" => rgb <= "101111";
					when "000111100100010" => rgb <= "101111";
					when "000111100100011" => rgb <= "101111";
					when "000111100100100" => rgb <= "101111";
					when "000111100100101" => rgb <= "001000";
					when "000111100100110" => rgb <= "001000";
					when "000111100100111" => rgb <= "001000";
					when "000111100101000" => rgb <= "000000";
					when "000111100101001" => rgb <= "000000";
					when "000111100101010" => rgb <= "000000";
					when "000111100101011" => rgb <= "000000";
					when "000111100101100" => rgb <= "000000";
					when "000111100101101" => rgb <= "000000";
					when "000111100101110" => rgb <= "000000";
					when "000111100101111" => rgb <= "000000";
					when "000111100110000" => rgb <= "000000";
					when "000111100110001" => rgb <= "000000";
					when "000111100110010" => rgb <= "000000";
					when "000111100110011" => rgb <= "000000";
					when "000111100110100" => rgb <= "000000";
					when "000111100110101" => rgb <= "000000";
					when "000111100110110" => rgb <= "000000";
					when "000111100110111" => rgb <= "000000";
					when "000111100111000" => rgb <= "000000";
					when "000111100111001" => rgb <= "000000";
					when "000111100111010" => rgb <= "000000";
					when "000111100111011" => rgb <= "000000";
					when "000111100111100" => rgb <= "000000";
					when "000111100111101" => rgb <= "000000";
					when "000111100111110" => rgb <= "000000";
					when "000111100111111" => rgb <= "000000";
					when "000111101000000" => rgb <= "000000";
					when "000111101000001" => rgb <= "000000";
					when "000111101000010" => rgb <= "000000";
					when "000111101000011" => rgb <= "000000";
					when "000111101000100" => rgb <= "000000";
					when "000111101000101" => rgb <= "000000";
					when "000111101000110" => rgb <= "000000";
					when "000111101000111" => rgb <= "000000";
					when "000111101001000" => rgb <= "000000";
					when "000111101001001" => rgb <= "000000";
					when "000111101001010" => rgb <= "000000";
					when "000111101001011" => rgb <= "000000";
					when "000111101001100" => rgb <= "000000";
					when "000111101001101" => rgb <= "000000";
					when "000111101001110" => rgb <= "000000";
					when "000111101001111" => rgb <= "000000";
					when "000111101010000" => rgb <= "000000";
					when "000111101010001" => rgb <= "000000";
					when "000111101010010" => rgb <= "000000";
					when "000111101010011" => rgb <= "000000";
					when "000111101010100" => rgb <= "000000";
					when "000111101010101" => rgb <= "000000";
					when "000111101010110" => rgb <= "000000";
					when "000111101010111" => rgb <= "000000";
					when "000111101011000" => rgb <= "000000";
					when "000111101011001" => rgb <= "000000";
					when "000111101011010" => rgb <= "000000";
					when "000111101011011" => rgb <= "000000";
					when "000111101011100" => rgb <= "000000";
					when "000111101011101" => rgb <= "000000";
					when "000111101011110" => rgb <= "000000";
					when "000111101011111" => rgb <= "000000";
					when "000111101100000" => rgb <= "000000";
					when "000111101100001" => rgb <= "000000";
					when "000111101100010" => rgb <= "000000";
					when "000111101100011" => rgb <= "000000";
					when "000111101100100" => rgb <= "000000";
					when "000111101100101" => rgb <= "000000";
					when "000111101100110" => rgb <= "000000";
					when "000111101100111" => rgb <= "000000";
					when "000111101101000" => rgb <= "000000";
					when "000111101101001" => rgb <= "000000";
					when "000111101101010" => rgb <= "000000";
					when "000111101101011" => rgb <= "000000";
					when "000111101101100" => rgb <= "000000";
					when "000111101101101" => rgb <= "000000";
					when "000111101101110" => rgb <= "000000";
					when "000111101101111" => rgb <= "000000";
					when "000111101110000" => rgb <= "000000";
					when "000111101110001" => rgb <= "000000";
					when "000111101110010" => rgb <= "000000";
					when "000111101110011" => rgb <= "000000";
					when "000111101110100" => rgb <= "000000";
					when "000111101110101" => rgb <= "000000";
					when "000111101110110" => rgb <= "000000";
					when "000111101110111" => rgb <= "000000";
					when "000111101111000" => rgb <= "101111";
					when "000111101111001" => rgb <= "101111";
					when "000111101111010" => rgb <= "101111";
					when "000111101111011" => rgb <= "101111";
					when "000111101111100" => rgb <= "101111";
					when "000111101111101" => rgb <= "101111";
					when "000111101111110" => rgb <= "101111";
					when "000111101111111" => rgb <= "101111";
					when "000111110000000" => rgb <= "101111";
					when "000111110000001" => rgb <= "101111";
					when "000111110000010" => rgb <= "101111";
					when "000111110000011" => rgb <= "101111";
					when "000111110000100" => rgb <= "101111";
					when "000111110000101" => rgb <= "101111";
					when "000111110000110" => rgb <= "101111";
					when "000111110000111" => rgb <= "101111";
					when "000111110001000" => rgb <= "101111";
					when "000111110001001" => rgb <= "101111";
					when "000111110001010" => rgb <= "101111";
					when "000111110001011" => rgb <= "101111";
					when "000111110001100" => rgb <= "101111";
					when "000111110001101" => rgb <= "101111";
					when "000111110001110" => rgb <= "101111";
					when "000111110001111" => rgb <= "101111";
					when "000111110010000" => rgb <= "101111";
					when "000111110010001" => rgb <= "101111";
					when "000111110010010" => rgb <= "101111";
					when "000111110010011" => rgb <= "101111";
					when "000111110010100" => rgb <= "101111";
					when "000111110010101" => rgb <= "101111";
					when "000111110010110" => rgb <= "101111";
					when "000111110010111" => rgb <= "101111";
					when "000111110011000" => rgb <= "101111";
					when "000111110011001" => rgb <= "101111";
					when "000111110011010" => rgb <= "101111";
					when "000111110011011" => rgb <= "101111";
					when "000111110011100" => rgb <= "101111";
					when "000111110011101" => rgb <= "101111";
					when "000111110011110" => rgb <= "101111";
					when "000111110011111" => rgb <= "101111";
					when "001000000000000" => rgb <= "101111";
					when "001000000000001" => rgb <= "101111";
					when "001000000000010" => rgb <= "000000";
					when "001000000000011" => rgb <= "000000";
					when "001000000000100" => rgb <= "001000";
					when "001000000000101" => rgb <= "001000";
					when "001000000000110" => rgb <= "001000";
					when "001000000000111" => rgb <= "001000";
					when "001000000001000" => rgb <= "001000";
					when "001000000001001" => rgb <= "001000";
					when "001000000001010" => rgb <= "001000";
					when "001000000001011" => rgb <= "001000";
					when "001000000001100" => rgb <= "001000";
					when "001000000001101" => rgb <= "001000";
					when "001000000001110" => rgb <= "001000";
					when "001000000001111" => rgb <= "001000";
					when "001000000010000" => rgb <= "001000";
					when "001000000010001" => rgb <= "001000";
					when "001000000010010" => rgb <= "001000";
					when "001000000010011" => rgb <= "001000";
					when "001000000010100" => rgb <= "001000";
					when "001000000010101" => rgb <= "001000";
					when "001000000010110" => rgb <= "001000";
					when "001000000010111" => rgb <= "001000";
					when "001000000011000" => rgb <= "001000";
					when "001000000011001" => rgb <= "001000";
					when "001000000011010" => rgb <= "001000";
					when "001000000011011" => rgb <= "001000";
					when "001000000011100" => rgb <= "001000";
					when "001000000011101" => rgb <= "001000";
					when "001000000011110" => rgb <= "001000";
					when "001000000011111" => rgb <= "001000";
					when "001000000100000" => rgb <= "001000";
					when "001000000100001" => rgb <= "001000";
					when "001000000100010" => rgb <= "001000";
					when "001000000100011" => rgb <= "001000";
					when "001000000100100" => rgb <= "001000";
					when "001000000100101" => rgb <= "001000";
					when "001000000100110" => rgb <= "001000";
					when "001000000100111" => rgb <= "001000";
					when "001000000101000" => rgb <= "001000";
					when "001000000101001" => rgb <= "001000";
					when "001000000101010" => rgb <= "001000";
					when "001000000101011" => rgb <= "001000";
					when "001000000101100" => rgb <= "001000";
					when "001000000101101" => rgb <= "001000";
					when "001000000101110" => rgb <= "001000";
					when "001000000101111" => rgb <= "001000";
					when "001000000110000" => rgb <= "001000";
					when "001000000110001" => rgb <= "001000";
					when "001000000110010" => rgb <= "001000";
					when "001000000110011" => rgb <= "001000";
					when "001000000110100" => rgb <= "001000";
					when "001000000110101" => rgb <= "001000";
					when "001000000110110" => rgb <= "001000";
					when "001000000110111" => rgb <= "001000";
					when "001000000111000" => rgb <= "001000";
					when "001000000111001" => rgb <= "001000";
					when "001000000111010" => rgb <= "001000";
					when "001000000111011" => rgb <= "001000";
					when "001000000111100" => rgb <= "001000";
					when "001000000111101" => rgb <= "001000";
					when "001000000111110" => rgb <= "001000";
					when "001000000111111" => rgb <= "001000";
					when "001000001000000" => rgb <= "001000";
					when "001000001000001" => rgb <= "001000";
					when "001000001000010" => rgb <= "001000";
					when "001000001000011" => rgb <= "001000";
					when "001000001000100" => rgb <= "001000";
					when "001000001000101" => rgb <= "001000";
					when "001000001000110" => rgb <= "001000";
					when "001000001000111" => rgb <= "001000";
					when "001000001001000" => rgb <= "001000";
					when "001000001001001" => rgb <= "001000";
					when "001000001001010" => rgb <= "000000";
					when "001000001001011" => rgb <= "000000";
					when "001000001001100" => rgb <= "000000";
					when "001000001001101" => rgb <= "000000";
					when "001000001001110" => rgb <= "101111";
					when "001000001001111" => rgb <= "101111";
					when "001000001010000" => rgb <= "101111";
					when "001000001010001" => rgb <= "101111";
					when "001000001010010" => rgb <= "101111";
					when "001000001010011" => rgb <= "101111";
					when "001000001010100" => rgb <= "101111";
					when "001000001010101" => rgb <= "101111";
					when "001000001010110" => rgb <= "101111";
					when "001000001010111" => rgb <= "101111";
					when "001000001011000" => rgb <= "101111";
					when "001000001011001" => rgb <= "101111";
					when "001000001011010" => rgb <= "101111";
					when "001000001011011" => rgb <= "101111";
					when "001000001011100" => rgb <= "101111";
					when "001000001011101" => rgb <= "101111";
					when "001000001011110" => rgb <= "101111";
					when "001000001011111" => rgb <= "101111";
					when "001000001100000" => rgb <= "101111";
					when "001000001100001" => rgb <= "101111";
					when "001000001100010" => rgb <= "101111";
					when "001000001100011" => rgb <= "101111";
					when "001000001100100" => rgb <= "101111";
					when "001000001100101" => rgb <= "101111";
					when "001000001100110" => rgb <= "101111";
					when "001000001100111" => rgb <= "101111";
					when "001000001101000" => rgb <= "101111";
					when "001000001101001" => rgb <= "101111";
					when "001000001101010" => rgb <= "101111";
					when "001000001101011" => rgb <= "101111";
					when "001000001101100" => rgb <= "101111";
					when "001000001101101" => rgb <= "101111";
					when "001000001101110" => rgb <= "101111";
					when "001000001101111" => rgb <= "101111";
					when "001000001110000" => rgb <= "101111";
					when "001000001110001" => rgb <= "101111";
					when "001000001110010" => rgb <= "101111";
					when "001000001110011" => rgb <= "101111";
					when "001000001110100" => rgb <= "101111";
					when "001000001110101" => rgb <= "101111";
					when "001000001110110" => rgb <= "101111";
					when "001000001110111" => rgb <= "101111";
					when "001000001111000" => rgb <= "101111";
					when "001000001111001" => rgb <= "101111";
					when "001000001111010" => rgb <= "101111";
					when "001000001111011" => rgb <= "101111";
					when "001000001111100" => rgb <= "101111";
					when "001000001111101" => rgb <= "101111";
					when "001000001111110" => rgb <= "101111";
					when "001000001111111" => rgb <= "101111";
					when "001000010000000" => rgb <= "101111";
					when "001000010000001" => rgb <= "101111";
					when "001000010000010" => rgb <= "101111";
					when "001000010000011" => rgb <= "101111";
					when "001000010000100" => rgb <= "101111";
					when "001000010000101" => rgb <= "101111";
					when "001000010000110" => rgb <= "101111";
					when "001000010000111" => rgb <= "101111";
					when "001000010001000" => rgb <= "101111";
					when "001000010001001" => rgb <= "101111";
					when "001000010001010" => rgb <= "101111";
					when "001000010001011" => rgb <= "101111";
					when "001000010001100" => rgb <= "101111";
					when "001000010001101" => rgb <= "101111";
					when "001000010001110" => rgb <= "101111";
					when "001000010001111" => rgb <= "101111";
					when "001000010010000" => rgb <= "101111";
					when "001000010010001" => rgb <= "101111";
					when "001000010010010" => rgb <= "101111";
					when "001000010010011" => rgb <= "101111";
					when "001000010010100" => rgb <= "101111";
					when "001000010010101" => rgb <= "101111";
					when "001000010010110" => rgb <= "101111";
					when "001000010010111" => rgb <= "101111";
					when "001000010011000" => rgb <= "101111";
					when "001000010011001" => rgb <= "101111";
					when "001000010011010" => rgb <= "101111";
					when "001000010011011" => rgb <= "101111";
					when "001000010011100" => rgb <= "101111";
					when "001000010011101" => rgb <= "101111";
					when "001000010011110" => rgb <= "101111";
					when "001000010011111" => rgb <= "101111";
					when "001000100000000" => rgb <= "101111";
					when "001000100000001" => rgb <= "101111";
					when "001000100000010" => rgb <= "000000";
					when "001000100000011" => rgb <= "000000";
					when "001000100000100" => rgb <= "001000";
					when "001000100000101" => rgb <= "001000";
					when "001000100000110" => rgb <= "001000";
					when "001000100000111" => rgb <= "001000";
					when "001000100001000" => rgb <= "001000";
					when "001000100001001" => rgb <= "001000";
					when "001000100001010" => rgb <= "001000";
					when "001000100001011" => rgb <= "001000";
					when "001000100001100" => rgb <= "001000";
					when "001000100001101" => rgb <= "001000";
					when "001000100001110" => rgb <= "001000";
					when "001000100001111" => rgb <= "001000";
					when "001000100010000" => rgb <= "001000";
					when "001000100010001" => rgb <= "001000";
					when "001000100010010" => rgb <= "001000";
					when "001000100010011" => rgb <= "001000";
					when "001000100010100" => rgb <= "001000";
					when "001000100010101" => rgb <= "001000";
					when "001000100010110" => rgb <= "001000";
					when "001000100010111" => rgb <= "001000";
					when "001000100011000" => rgb <= "001000";
					when "001000100011001" => rgb <= "001000";
					when "001000100011010" => rgb <= "001000";
					when "001000100011011" => rgb <= "001000";
					when "001000100011100" => rgb <= "001000";
					when "001000100011101" => rgb <= "001000";
					when "001000100011110" => rgb <= "001000";
					when "001000100011111" => rgb <= "001000";
					when "001000100100000" => rgb <= "001000";
					when "001000100100001" => rgb <= "001000";
					when "001000100100010" => rgb <= "001000";
					when "001000100100011" => rgb <= "001000";
					when "001000100100100" => rgb <= "001000";
					when "001000100100101" => rgb <= "001000";
					when "001000100100110" => rgb <= "001000";
					when "001000100100111" => rgb <= "001000";
					when "001000100101000" => rgb <= "001000";
					when "001000100101001" => rgb <= "001000";
					when "001000100101010" => rgb <= "001000";
					when "001000100101011" => rgb <= "001000";
					when "001000100101100" => rgb <= "001000";
					when "001000100101101" => rgb <= "001000";
					when "001000100101110" => rgb <= "001000";
					when "001000100101111" => rgb <= "001000";
					when "001000100110000" => rgb <= "001000";
					when "001000100110001" => rgb <= "001000";
					when "001000100110010" => rgb <= "001000";
					when "001000100110011" => rgb <= "001000";
					when "001000100110100" => rgb <= "001000";
					when "001000100110101" => rgb <= "001000";
					when "001000100110110" => rgb <= "001000";
					when "001000100110111" => rgb <= "001000";
					when "001000100111000" => rgb <= "001000";
					when "001000100111001" => rgb <= "001000";
					when "001000100111010" => rgb <= "001000";
					when "001000100111011" => rgb <= "001000";
					when "001000100111100" => rgb <= "001000";
					when "001000100111101" => rgb <= "001000";
					when "001000100111110" => rgb <= "001000";
					when "001000100111111" => rgb <= "001000";
					when "001000101000000" => rgb <= "001000";
					when "001000101000001" => rgb <= "001000";
					when "001000101000010" => rgb <= "001000";
					when "001000101000011" => rgb <= "001000";
					when "001000101000100" => rgb <= "001000";
					when "001000101000101" => rgb <= "001000";
					when "001000101000110" => rgb <= "001000";
					when "001000101000111" => rgb <= "001000";
					when "001000101001000" => rgb <= "001000";
					when "001000101001001" => rgb <= "001000";
					when "001000101001010" => rgb <= "000000";
					when "001000101001011" => rgb <= "000000";
					when "001000101001100" => rgb <= "000000";
					when "001000101001101" => rgb <= "000000";
					when "001000101001110" => rgb <= "101111";
					when "001000101001111" => rgb <= "101111";
					when "001000101010000" => rgb <= "101111";
					when "001000101010001" => rgb <= "101111";
					when "001000101010010" => rgb <= "101111";
					when "001000101010011" => rgb <= "101111";
					when "001000101010100" => rgb <= "101111";
					when "001000101010101" => rgb <= "101111";
					when "001000101010110" => rgb <= "101111";
					when "001000101010111" => rgb <= "101111";
					when "001000101011000" => rgb <= "101111";
					when "001000101011001" => rgb <= "101111";
					when "001000101011010" => rgb <= "101111";
					when "001000101011011" => rgb <= "101111";
					when "001000101011100" => rgb <= "101111";
					when "001000101011101" => rgb <= "101111";
					when "001000101011110" => rgb <= "101111";
					when "001000101011111" => rgb <= "101111";
					when "001000101100000" => rgb <= "101111";
					when "001000101100001" => rgb <= "101111";
					when "001000101100010" => rgb <= "101111";
					when "001000101100011" => rgb <= "101111";
					when "001000101100100" => rgb <= "101111";
					when "001000101100101" => rgb <= "101111";
					when "001000101100110" => rgb <= "101111";
					when "001000101100111" => rgb <= "101111";
					when "001000101101000" => rgb <= "101111";
					when "001000101101001" => rgb <= "101111";
					when "001000101101010" => rgb <= "101111";
					when "001000101101011" => rgb <= "101111";
					when "001000101101100" => rgb <= "101111";
					when "001000101101101" => rgb <= "101111";
					when "001000101101110" => rgb <= "101111";
					when "001000101101111" => rgb <= "101111";
					when "001000101110000" => rgb <= "101111";
					when "001000101110001" => rgb <= "101111";
					when "001000101110010" => rgb <= "101111";
					when "001000101110011" => rgb <= "101111";
					when "001000101110100" => rgb <= "101111";
					when "001000101110101" => rgb <= "101111";
					when "001000101110110" => rgb <= "101111";
					when "001000101110111" => rgb <= "101111";
					when "001000101111000" => rgb <= "101111";
					when "001000101111001" => rgb <= "101111";
					when "001000101111010" => rgb <= "101111";
					when "001000101111011" => rgb <= "101111";
					when "001000101111100" => rgb <= "101111";
					when "001000101111101" => rgb <= "101111";
					when "001000101111110" => rgb <= "101111";
					when "001000101111111" => rgb <= "101111";
					when "001000110000000" => rgb <= "101111";
					when "001000110000001" => rgb <= "101111";
					when "001000110000010" => rgb <= "101111";
					when "001000110000011" => rgb <= "101111";
					when "001000110000100" => rgb <= "101111";
					when "001000110000101" => rgb <= "101111";
					when "001000110000110" => rgb <= "101111";
					when "001000110000111" => rgb <= "101111";
					when "001000110001000" => rgb <= "101111";
					when "001000110001001" => rgb <= "101111";
					when "001000110001010" => rgb <= "101111";
					when "001000110001011" => rgb <= "101111";
					when "001000110001100" => rgb <= "101111";
					when "001000110001101" => rgb <= "101111";
					when "001000110001110" => rgb <= "101111";
					when "001000110001111" => rgb <= "101111";
					when "001000110010000" => rgb <= "101111";
					when "001000110010001" => rgb <= "101111";
					when "001000110010010" => rgb <= "101111";
					when "001000110010011" => rgb <= "101111";
					when "001000110010100" => rgb <= "101111";
					when "001000110010101" => rgb <= "101111";
					when "001000110010110" => rgb <= "101111";
					when "001000110010111" => rgb <= "101111";
					when "001000110011000" => rgb <= "101111";
					when "001000110011001" => rgb <= "101111";
					when "001000110011010" => rgb <= "101111";
					when "001000110011011" => rgb <= "101111";
					when "001000110011100" => rgb <= "101111";
					when "001000110011101" => rgb <= "101111";
					when "001000110011110" => rgb <= "101111";
					when "001000110011111" => rgb <= "101111";
					when "001001000000000" => rgb <= "000000";
					when "001001000000001" => rgb <= "000000";
					when "001001000000010" => rgb <= "000000";
					when "001001000000011" => rgb <= "000000";
					when "001001000000100" => rgb <= "001000";
					when "001001000000101" => rgb <= "001000";
					when "001001000000110" => rgb <= "001000";
					when "001001000000111" => rgb <= "001000";
					when "001001000001000" => rgb <= "001000";
					when "001001000001001" => rgb <= "001000";
					when "001001000001010" => rgb <= "001000";
					when "001001000001011" => rgb <= "001000";
					when "001001000001100" => rgb <= "001000";
					when "001001000001101" => rgb <= "001000";
					when "001001000001110" => rgb <= "001000";
					when "001001000001111" => rgb <= "001000";
					when "001001000010000" => rgb <= "001000";
					when "001001000010001" => rgb <= "001000";
					when "001001000010010" => rgb <= "001000";
					when "001001000010011" => rgb <= "001000";
					when "001001000010100" => rgb <= "001000";
					when "001001000010101" => rgb <= "001000";
					when "001001000010110" => rgb <= "001000";
					when "001001000010111" => rgb <= "001000";
					when "001001000011000" => rgb <= "001000";
					when "001001000011001" => rgb <= "001000";
					when "001001000011010" => rgb <= "001000";
					when "001001000011011" => rgb <= "001000";
					when "001001000011100" => rgb <= "001000";
					when "001001000011101" => rgb <= "001000";
					when "001001000011110" => rgb <= "001000";
					when "001001000011111" => rgb <= "001000";
					when "001001000100000" => rgb <= "001000";
					when "001001000100001" => rgb <= "001000";
					when "001001000100010" => rgb <= "001000";
					when "001001000100011" => rgb <= "001000";
					when "001001000100100" => rgb <= "001000";
					when "001001000100101" => rgb <= "001000";
					when "001001000100110" => rgb <= "001000";
					when "001001000100111" => rgb <= "001000";
					when "001001000101000" => rgb <= "001000";
					when "001001000101001" => rgb <= "001000";
					when "001001000101010" => rgb <= "001000";
					when "001001000101011" => rgb <= "001000";
					when "001001000101100" => rgb <= "001000";
					when "001001000101101" => rgb <= "001000";
					when "001001000101110" => rgb <= "001000";
					when "001001000101111" => rgb <= "001000";
					when "001001000110000" => rgb <= "001000";
					when "001001000110001" => rgb <= "001000";
					when "001001000110010" => rgb <= "001000";
					when "001001000110011" => rgb <= "001000";
					when "001001000110100" => rgb <= "001000";
					when "001001000110101" => rgb <= "001000";
					when "001001000110110" => rgb <= "001000";
					when "001001000110111" => rgb <= "001000";
					when "001001000111000" => rgb <= "001000";
					when "001001000111001" => rgb <= "001000";
					when "001001000111010" => rgb <= "001000";
					when "001001000111011" => rgb <= "001000";
					when "001001000111100" => rgb <= "001000";
					when "001001000111101" => rgb <= "001000";
					when "001001000111110" => rgb <= "001000";
					when "001001000111111" => rgb <= "001000";
					when "001001001000000" => rgb <= "001000";
					when "001001001000001" => rgb <= "001000";
					when "001001001000010" => rgb <= "001000";
					when "001001001000011" => rgb <= "001000";
					when "001001001000100" => rgb <= "001000";
					when "001001001000101" => rgb <= "001000";
					when "001001001000110" => rgb <= "001000";
					when "001001001000111" => rgb <= "001000";
					when "001001001001000" => rgb <= "001000";
					when "001001001001001" => rgb <= "001000";
					when "001001001001010" => rgb <= "001000";
					when "001001001001011" => rgb <= "001000";
					when "001001001001100" => rgb <= "001000";
					when "001001001001101" => rgb <= "001000";
					when "001001001001110" => rgb <= "000000";
					when "001001001001111" => rgb <= "000000";
					when "001001001010000" => rgb <= "101111";
					when "001001001010001" => rgb <= "101111";
					when "001001001010010" => rgb <= "101111";
					when "001001001010011" => rgb <= "101111";
					when "001001001010100" => rgb <= "101111";
					when "001001001010101" => rgb <= "101111";
					when "001001001010110" => rgb <= "101111";
					when "001001001010111" => rgb <= "101111";
					when "001001001011000" => rgb <= "101111";
					when "001001001011001" => rgb <= "101111";
					when "001001001011010" => rgb <= "101111";
					when "001001001011011" => rgb <= "101111";
					when "001001001011100" => rgb <= "101111";
					when "001001001011101" => rgb <= "101111";
					when "001001001011110" => rgb <= "101111";
					when "001001001011111" => rgb <= "101111";
					when "001001001100000" => rgb <= "101111";
					when "001001001100001" => rgb <= "101111";
					when "001001001100010" => rgb <= "101111";
					when "001001001100011" => rgb <= "101111";
					when "001001001100100" => rgb <= "101111";
					when "001001001100101" => rgb <= "101111";
					when "001001001100110" => rgb <= "101111";
					when "001001001100111" => rgb <= "101111";
					when "001001001101000" => rgb <= "101111";
					when "001001001101001" => rgb <= "101111";
					when "001001001101010" => rgb <= "101111";
					when "001001001101011" => rgb <= "101111";
					when "001001001101100" => rgb <= "101111";
					when "001001001101101" => rgb <= "101111";
					when "001001001101110" => rgb <= "101111";
					when "001001001101111" => rgb <= "101111";
					when "001001001110000" => rgb <= "101111";
					when "001001001110001" => rgb <= "101111";
					when "001001001110010" => rgb <= "101111";
					when "001001001110011" => rgb <= "101111";
					when "001001001110100" => rgb <= "101111";
					when "001001001110101" => rgb <= "101111";
					when "001001001110110" => rgb <= "101111";
					when "001001001110111" => rgb <= "101111";
					when "001001001111000" => rgb <= "101111";
					when "001001001111001" => rgb <= "101111";
					when "001001001111010" => rgb <= "101111";
					when "001001001111011" => rgb <= "101111";
					when "001001001111100" => rgb <= "101111";
					when "001001001111101" => rgb <= "101111";
					when "001001001111110" => rgb <= "101111";
					when "001001001111111" => rgb <= "101111";
					when "001001010000000" => rgb <= "101111";
					when "001001010000001" => rgb <= "101111";
					when "001001010000010" => rgb <= "101111";
					when "001001010000011" => rgb <= "101111";
					when "001001010000100" => rgb <= "101111";
					when "001001010000101" => rgb <= "101111";
					when "001001010000110" => rgb <= "101111";
					when "001001010000111" => rgb <= "101111";
					when "001001010001000" => rgb <= "101111";
					when "001001010001001" => rgb <= "101111";
					when "001001010001010" => rgb <= "101111";
					when "001001010001011" => rgb <= "101111";
					when "001001010001100" => rgb <= "101111";
					when "001001010001101" => rgb <= "101111";
					when "001001010001110" => rgb <= "101111";
					when "001001010001111" => rgb <= "101111";
					when "001001010010000" => rgb <= "101111";
					when "001001010010001" => rgb <= "101111";
					when "001001010010010" => rgb <= "101111";
					when "001001010010011" => rgb <= "101111";
					when "001001010010100" => rgb <= "101111";
					when "001001010010101" => rgb <= "101111";
					when "001001010010110" => rgb <= "101111";
					when "001001010010111" => rgb <= "101111";
					when "001001010011000" => rgb <= "101111";
					when "001001010011001" => rgb <= "101111";
					when "001001010011010" => rgb <= "101111";
					when "001001010011011" => rgb <= "101111";
					when "001001010011100" => rgb <= "101111";
					when "001001010011101" => rgb <= "101111";
					when "001001010011110" => rgb <= "101111";
					when "001001010011111" => rgb <= "101111";
					when "001001100000000" => rgb <= "000000";
					when "001001100000001" => rgb <= "000000";
					when "001001100000010" => rgb <= "000000";
					when "001001100000011" => rgb <= "000000";
					when "001001100000100" => rgb <= "001000";
					when "001001100000101" => rgb <= "001000";
					when "001001100000110" => rgb <= "001000";
					when "001001100000111" => rgb <= "001000";
					when "001001100001000" => rgb <= "001000";
					when "001001100001001" => rgb <= "001000";
					when "001001100001010" => rgb <= "001000";
					when "001001100001011" => rgb <= "001000";
					when "001001100001100" => rgb <= "001000";
					when "001001100001101" => rgb <= "001000";
					when "001001100001110" => rgb <= "001000";
					when "001001100001111" => rgb <= "001000";
					when "001001100010000" => rgb <= "001000";
					when "001001100010001" => rgb <= "001000";
					when "001001100010010" => rgb <= "001000";
					when "001001100010011" => rgb <= "001000";
					when "001001100010100" => rgb <= "001000";
					when "001001100010101" => rgb <= "001000";
					when "001001100010110" => rgb <= "001000";
					when "001001100010111" => rgb <= "001000";
					when "001001100011000" => rgb <= "001000";
					when "001001100011001" => rgb <= "001000";
					when "001001100011010" => rgb <= "001000";
					when "001001100011011" => rgb <= "001000";
					when "001001100011100" => rgb <= "001000";
					when "001001100011101" => rgb <= "001000";
					when "001001100011110" => rgb <= "001000";
					when "001001100011111" => rgb <= "001000";
					when "001001100100000" => rgb <= "001000";
					when "001001100100001" => rgb <= "001000";
					when "001001100100010" => rgb <= "001000";
					when "001001100100011" => rgb <= "001000";
					when "001001100100100" => rgb <= "001000";
					when "001001100100101" => rgb <= "001000";
					when "001001100100110" => rgb <= "001000";
					when "001001100100111" => rgb <= "001000";
					when "001001100101000" => rgb <= "001000";
					when "001001100101001" => rgb <= "001000";
					when "001001100101010" => rgb <= "001000";
					when "001001100101011" => rgb <= "001000";
					when "001001100101100" => rgb <= "001000";
					when "001001100101101" => rgb <= "001000";
					when "001001100101110" => rgb <= "001000";
					when "001001100101111" => rgb <= "001000";
					when "001001100110000" => rgb <= "001000";
					when "001001100110001" => rgb <= "001000";
					when "001001100110010" => rgb <= "001000";
					when "001001100110011" => rgb <= "001000";
					when "001001100110100" => rgb <= "001000";
					when "001001100110101" => rgb <= "001000";
					when "001001100110110" => rgb <= "001000";
					when "001001100110111" => rgb <= "001000";
					when "001001100111000" => rgb <= "001000";
					when "001001100111001" => rgb <= "001000";
					when "001001100111010" => rgb <= "001000";
					when "001001100111011" => rgb <= "001000";
					when "001001100111100" => rgb <= "001000";
					when "001001100111101" => rgb <= "001000";
					when "001001100111110" => rgb <= "001000";
					when "001001100111111" => rgb <= "001000";
					when "001001101000000" => rgb <= "001000";
					when "001001101000001" => rgb <= "001000";
					when "001001101000010" => rgb <= "001000";
					when "001001101000011" => rgb <= "001000";
					when "001001101000100" => rgb <= "001000";
					when "001001101000101" => rgb <= "001000";
					when "001001101000110" => rgb <= "001000";
					when "001001101000111" => rgb <= "001000";
					when "001001101001000" => rgb <= "001000";
					when "001001101001001" => rgb <= "001000";
					when "001001101001010" => rgb <= "001000";
					when "001001101001011" => rgb <= "001000";
					when "001001101001100" => rgb <= "001000";
					when "001001101001101" => rgb <= "001000";
					when "001001101001110" => rgb <= "000000";
					when "001001101001111" => rgb <= "000000";
					when "001001101010000" => rgb <= "101111";
					when "001001101010001" => rgb <= "101111";
					when "001001101010010" => rgb <= "101111";
					when "001001101010011" => rgb <= "101111";
					when "001001101010100" => rgb <= "101111";
					when "001001101010101" => rgb <= "101111";
					when "001001101010110" => rgb <= "101111";
					when "001001101010111" => rgb <= "101111";
					when "001001101011000" => rgb <= "101111";
					when "001001101011001" => rgb <= "101111";
					when "001001101011010" => rgb <= "101111";
					when "001001101011011" => rgb <= "101111";
					when "001001101011100" => rgb <= "101111";
					when "001001101011101" => rgb <= "101111";
					when "001001101011110" => rgb <= "101111";
					when "001001101011111" => rgb <= "101111";
					when "001001101100000" => rgb <= "101111";
					when "001001101100001" => rgb <= "101111";
					when "001001101100010" => rgb <= "101111";
					when "001001101100011" => rgb <= "101111";
					when "001001101100100" => rgb <= "101111";
					when "001001101100101" => rgb <= "101111";
					when "001001101100110" => rgb <= "101111";
					when "001001101100111" => rgb <= "101111";
					when "001001101101000" => rgb <= "101111";
					when "001001101101001" => rgb <= "101111";
					when "001001101101010" => rgb <= "101111";
					when "001001101101011" => rgb <= "101111";
					when "001001101101100" => rgb <= "101111";
					when "001001101101101" => rgb <= "101111";
					when "001001101101110" => rgb <= "101111";
					when "001001101101111" => rgb <= "101111";
					when "001001101110000" => rgb <= "101111";
					when "001001101110001" => rgb <= "101111";
					when "001001101110010" => rgb <= "101111";
					when "001001101110011" => rgb <= "101111";
					when "001001101110100" => rgb <= "101111";
					when "001001101110101" => rgb <= "101111";
					when "001001101110110" => rgb <= "101111";
					when "001001101110111" => rgb <= "101111";
					when "001001101111000" => rgb <= "101111";
					when "001001101111001" => rgb <= "101111";
					when "001001101111010" => rgb <= "101111";
					when "001001101111011" => rgb <= "101111";
					when "001001101111100" => rgb <= "101111";
					when "001001101111101" => rgb <= "101111";
					when "001001101111110" => rgb <= "101111";
					when "001001101111111" => rgb <= "101111";
					when "001001110000000" => rgb <= "101111";
					when "001001110000001" => rgb <= "101111";
					when "001001110000010" => rgb <= "101111";
					when "001001110000011" => rgb <= "101111";
					when "001001110000100" => rgb <= "101111";
					when "001001110000101" => rgb <= "101111";
					when "001001110000110" => rgb <= "101111";
					when "001001110000111" => rgb <= "101111";
					when "001001110001000" => rgb <= "101111";
					when "001001110001001" => rgb <= "101111";
					when "001001110001010" => rgb <= "101111";
					when "001001110001011" => rgb <= "101111";
					when "001001110001100" => rgb <= "101111";
					when "001001110001101" => rgb <= "101111";
					when "001001110001110" => rgb <= "101111";
					when "001001110001111" => rgb <= "101111";
					when "001001110010000" => rgb <= "101111";
					when "001001110010001" => rgb <= "101111";
					when "001001110010010" => rgb <= "101111";
					when "001001110010011" => rgb <= "101111";
					when "001001110010100" => rgb <= "101111";
					when "001001110010101" => rgb <= "101111";
					when "001001110010110" => rgb <= "101111";
					when "001001110010111" => rgb <= "101111";
					when "001001110011000" => rgb <= "101111";
					when "001001110011001" => rgb <= "101111";
					when "001001110011010" => rgb <= "101111";
					when "001001110011011" => rgb <= "101111";
					when "001001110011100" => rgb <= "101111";
					when "001001110011101" => rgb <= "101111";
					when "001001110011110" => rgb <= "101111";
					when "001001110011111" => rgb <= "101111";
					when "001010000000000" => rgb <= "001000";
					when "001010000000001" => rgb <= "001000";
					when "001010000000010" => rgb <= "001000";
					when "001010000000011" => rgb <= "001000";
					when "001010000000100" => rgb <= "001000";
					when "001010000000101" => rgb <= "001000";
					when "001010000000110" => rgb <= "001000";
					when "001010000000111" => rgb <= "001000";
					when "001010000001000" => rgb <= "001000";
					when "001010000001001" => rgb <= "001000";
					when "001010000001010" => rgb <= "001000";
					when "001010000001011" => rgb <= "001000";
					when "001010000001100" => rgb <= "001000";
					when "001010000001101" => rgb <= "001000";
					when "001010000001110" => rgb <= "001000";
					when "001010000001111" => rgb <= "001000";
					when "001010000010000" => rgb <= "001000";
					when "001010000010001" => rgb <= "001000";
					when "001010000010010" => rgb <= "001000";
					when "001010000010011" => rgb <= "001000";
					when "001010000010100" => rgb <= "001000";
					when "001010000010101" => rgb <= "001000";
					when "001010000010110" => rgb <= "001000";
					when "001010000010111" => rgb <= "001000";
					when "001010000011000" => rgb <= "001000";
					when "001010000011001" => rgb <= "001000";
					when "001010000011010" => rgb <= "001000";
					when "001010000011011" => rgb <= "001000";
					when "001010000011100" => rgb <= "001000";
					when "001010000011101" => rgb <= "001000";
					when "001010000011110" => rgb <= "001000";
					when "001010000011111" => rgb <= "001000";
					when "001010000100000" => rgb <= "001000";
					when "001010000100001" => rgb <= "001000";
					when "001010000100010" => rgb <= "001000";
					when "001010000100011" => rgb <= "001000";
					when "001010000100100" => rgb <= "001000";
					when "001010000100101" => rgb <= "001000";
					when "001010000100110" => rgb <= "001000";
					when "001010000100111" => rgb <= "001000";
					when "001010000101000" => rgb <= "001000";
					when "001010000101001" => rgb <= "001000";
					when "001010000101010" => rgb <= "001000";
					when "001010000101011" => rgb <= "001000";
					when "001010000101100" => rgb <= "001000";
					when "001010000101101" => rgb <= "001000";
					when "001010000101110" => rgb <= "001000";
					when "001010000101111" => rgb <= "001000";
					when "001010000110000" => rgb <= "001000";
					when "001010000110001" => rgb <= "001000";
					when "001010000110010" => rgb <= "001000";
					when "001010000110011" => rgb <= "001000";
					when "001010000110100" => rgb <= "001000";
					when "001010000110101" => rgb <= "001000";
					when "001010000110110" => rgb <= "001000";
					when "001010000110111" => rgb <= "001000";
					when "001010000111000" => rgb <= "001000";
					when "001010000111001" => rgb <= "001000";
					when "001010000111010" => rgb <= "001000";
					when "001010000111011" => rgb <= "001000";
					when "001010000111100" => rgb <= "001000";
					when "001010000111101" => rgb <= "001000";
					when "001010000111110" => rgb <= "001000";
					when "001010000111111" => rgb <= "001000";
					when "001010001000000" => rgb <= "001000";
					when "001010001000001" => rgb <= "001000";
					when "001010001000010" => rgb <= "001000";
					when "001010001000011" => rgb <= "001000";
					when "001010001000100" => rgb <= "001000";
					when "001010001000101" => rgb <= "001000";
					when "001010001000110" => rgb <= "001000";
					when "001010001000111" => rgb <= "001000";
					when "001010001001000" => rgb <= "001000";
					when "001010001001001" => rgb <= "001000";
					when "001010001001010" => rgb <= "001000";
					when "001010001001011" => rgb <= "001000";
					when "001010001001100" => rgb <= "001000";
					when "001010001001101" => rgb <= "001000";
					when "001010001001110" => rgb <= "001000";
					when "001010001001111" => rgb <= "001000";
					when "001010001010000" => rgb <= "000000";
					when "001010001010001" => rgb <= "000000";
					when "001010001010010" => rgb <= "101111";
					when "001010001010011" => rgb <= "101111";
					when "001010001010100" => rgb <= "101111";
					when "001010001010101" => rgb <= "101111";
					when "001010001010110" => rgb <= "101111";
					when "001010001010111" => rgb <= "101111";
					when "001010001011000" => rgb <= "101111";
					when "001010001011001" => rgb <= "101111";
					when "001010001011010" => rgb <= "101111";
					when "001010001011011" => rgb <= "101111";
					when "001010001011100" => rgb <= "101111";
					when "001010001011101" => rgb <= "101111";
					when "001010001011110" => rgb <= "101111";
					when "001010001011111" => rgb <= "101111";
					when "001010001100000" => rgb <= "101111";
					when "001010001100001" => rgb <= "101111";
					when "001010001100010" => rgb <= "101111";
					when "001010001100011" => rgb <= "101111";
					when "001010001100100" => rgb <= "101111";
					when "001010001100101" => rgb <= "101111";
					when "001010001100110" => rgb <= "101111";
					when "001010001100111" => rgb <= "101111";
					when "001010001101000" => rgb <= "101111";
					when "001010001101001" => rgb <= "101111";
					when "001010001101010" => rgb <= "101111";
					when "001010001101011" => rgb <= "101111";
					when "001010001101100" => rgb <= "101111";
					when "001010001101101" => rgb <= "101111";
					when "001010001101110" => rgb <= "101111";
					when "001010001101111" => rgb <= "101111";
					when "001010001110000" => rgb <= "101111";
					when "001010001110001" => rgb <= "101111";
					when "001010001110010" => rgb <= "101111";
					when "001010001110011" => rgb <= "101111";
					when "001010001110100" => rgb <= "101111";
					when "001010001110101" => rgb <= "101111";
					when "001010001110110" => rgb <= "101111";
					when "001010001110111" => rgb <= "101111";
					when "001010001111000" => rgb <= "101111";
					when "001010001111001" => rgb <= "101111";
					when "001010001111010" => rgb <= "101111";
					when "001010001111011" => rgb <= "101111";
					when "001010001111100" => rgb <= "101111";
					when "001010001111101" => rgb <= "101111";
					when "001010001111110" => rgb <= "101111";
					when "001010001111111" => rgb <= "101111";
					when "001010010000000" => rgb <= "101111";
					when "001010010000001" => rgb <= "101111";
					when "001010010000010" => rgb <= "101111";
					when "001010010000011" => rgb <= "101111";
					when "001010010000100" => rgb <= "101111";
					when "001010010000101" => rgb <= "101111";
					when "001010010000110" => rgb <= "101111";
					when "001010010000111" => rgb <= "101111";
					when "001010010001000" => rgb <= "101111";
					when "001010010001001" => rgb <= "101111";
					when "001010010001010" => rgb <= "101111";
					when "001010010001011" => rgb <= "101111";
					when "001010010001100" => rgb <= "101111";
					when "001010010001101" => rgb <= "101111";
					when "001010010001110" => rgb <= "101111";
					when "001010010001111" => rgb <= "101111";
					when "001010010010000" => rgb <= "101111";
					when "001010010010001" => rgb <= "101111";
					when "001010010010010" => rgb <= "101111";
					when "001010010010011" => rgb <= "101111";
					when "001010010010100" => rgb <= "101111";
					when "001010010010101" => rgb <= "101111";
					when "001010010010110" => rgb <= "101111";
					when "001010010010111" => rgb <= "101111";
					when "001010010011000" => rgb <= "101111";
					when "001010010011001" => rgb <= "101111";
					when "001010010011010" => rgb <= "101111";
					when "001010010011011" => rgb <= "101111";
					when "001010010011100" => rgb <= "101111";
					when "001010010011101" => rgb <= "101111";
					when "001010010011110" => rgb <= "101111";
					when "001010010011111" => rgb <= "101111";
					when "001010100000000" => rgb <= "001000";
					when "001010100000001" => rgb <= "001000";
					when "001010100000010" => rgb <= "001000";
					when "001010100000011" => rgb <= "001000";
					when "001010100000100" => rgb <= "001000";
					when "001010100000101" => rgb <= "001000";
					when "001010100000110" => rgb <= "001000";
					when "001010100000111" => rgb <= "001000";
					when "001010100001000" => rgb <= "001000";
					when "001010100001001" => rgb <= "001000";
					when "001010100001010" => rgb <= "001000";
					when "001010100001011" => rgb <= "001000";
					when "001010100001100" => rgb <= "001000";
					when "001010100001101" => rgb <= "001000";
					when "001010100001110" => rgb <= "001000";
					when "001010100001111" => rgb <= "001000";
					when "001010100010000" => rgb <= "001000";
					when "001010100010001" => rgb <= "001000";
					when "001010100010010" => rgb <= "001000";
					when "001010100010011" => rgb <= "001000";
					when "001010100010100" => rgb <= "001000";
					when "001010100010101" => rgb <= "001000";
					when "001010100010110" => rgb <= "001000";
					when "001010100010111" => rgb <= "001000";
					when "001010100011000" => rgb <= "001000";
					when "001010100011001" => rgb <= "001000";
					when "001010100011010" => rgb <= "001000";
					when "001010100011011" => rgb <= "001000";
					when "001010100011100" => rgb <= "001000";
					when "001010100011101" => rgb <= "001000";
					when "001010100011110" => rgb <= "001000";
					when "001010100011111" => rgb <= "001000";
					when "001010100100000" => rgb <= "001000";
					when "001010100100001" => rgb <= "001000";
					when "001010100100010" => rgb <= "001000";
					when "001010100100011" => rgb <= "001000";
					when "001010100100100" => rgb <= "001000";
					when "001010100100101" => rgb <= "001000";
					when "001010100100110" => rgb <= "001000";
					when "001010100100111" => rgb <= "001000";
					when "001010100101000" => rgb <= "001000";
					when "001010100101001" => rgb <= "001000";
					when "001010100101010" => rgb <= "001000";
					when "001010100101011" => rgb <= "001000";
					when "001010100101100" => rgb <= "001000";
					when "001010100101101" => rgb <= "001000";
					when "001010100101110" => rgb <= "001000";
					when "001010100101111" => rgb <= "001000";
					when "001010100110000" => rgb <= "001000";
					when "001010100110001" => rgb <= "001000";
					when "001010100110010" => rgb <= "001000";
					when "001010100110011" => rgb <= "001000";
					when "001010100110100" => rgb <= "001000";
					when "001010100110101" => rgb <= "001000";
					when "001010100110110" => rgb <= "001000";
					when "001010100110111" => rgb <= "001000";
					when "001010100111000" => rgb <= "001000";
					when "001010100111001" => rgb <= "001000";
					when "001010100111010" => rgb <= "001000";
					when "001010100111011" => rgb <= "001000";
					when "001010100111100" => rgb <= "001000";
					when "001010100111101" => rgb <= "001000";
					when "001010100111110" => rgb <= "001000";
					when "001010100111111" => rgb <= "001000";
					when "001010101000000" => rgb <= "001000";
					when "001010101000001" => rgb <= "001000";
					when "001010101000010" => rgb <= "001000";
					when "001010101000011" => rgb <= "001000";
					when "001010101000100" => rgb <= "001000";
					when "001010101000101" => rgb <= "001000";
					when "001010101000110" => rgb <= "001000";
					when "001010101000111" => rgb <= "001000";
					when "001010101001000" => rgb <= "001000";
					when "001010101001001" => rgb <= "001000";
					when "001010101001010" => rgb <= "001000";
					when "001010101001011" => rgb <= "001000";
					when "001010101001100" => rgb <= "001000";
					when "001010101001101" => rgb <= "001000";
					when "001010101001110" => rgb <= "001000";
					when "001010101001111" => rgb <= "001000";
					when "001010101010000" => rgb <= "000000";
					when "001010101010001" => rgb <= "000000";
					when "001010101010010" => rgb <= "101111";
					when "001010101010011" => rgb <= "101111";
					when "001010101010100" => rgb <= "101111";
					when "001010101010101" => rgb <= "101111";
					when "001010101010110" => rgb <= "101111";
					when "001010101010111" => rgb <= "101111";
					when "001010101011000" => rgb <= "101111";
					when "001010101011001" => rgb <= "101111";
					when "001010101011010" => rgb <= "101111";
					when "001010101011011" => rgb <= "101111";
					when "001010101011100" => rgb <= "101111";
					when "001010101011101" => rgb <= "101111";
					when "001010101011110" => rgb <= "101111";
					when "001010101011111" => rgb <= "101111";
					when "001010101100000" => rgb <= "101111";
					when "001010101100001" => rgb <= "101111";
					when "001010101100010" => rgb <= "101111";
					when "001010101100011" => rgb <= "101111";
					when "001010101100100" => rgb <= "101111";
					when "001010101100101" => rgb <= "101111";
					when "001010101100110" => rgb <= "101111";
					when "001010101100111" => rgb <= "101111";
					when "001010101101000" => rgb <= "101111";
					when "001010101101001" => rgb <= "101111";
					when "001010101101010" => rgb <= "101111";
					when "001010101101011" => rgb <= "101111";
					when "001010101101100" => rgb <= "101111";
					when "001010101101101" => rgb <= "101111";
					when "001010101101110" => rgb <= "101111";
					when "001010101101111" => rgb <= "101111";
					when "001010101110000" => rgb <= "101111";
					when "001010101110001" => rgb <= "101111";
					when "001010101110010" => rgb <= "101111";
					when "001010101110011" => rgb <= "101111";
					when "001010101110100" => rgb <= "101111";
					when "001010101110101" => rgb <= "101111";
					when "001010101110110" => rgb <= "101111";
					when "001010101110111" => rgb <= "101111";
					when "001010101111000" => rgb <= "101111";
					when "001010101111001" => rgb <= "101111";
					when "001010101111010" => rgb <= "101111";
					when "001010101111011" => rgb <= "101111";
					when "001010101111100" => rgb <= "101111";
					when "001010101111101" => rgb <= "101111";
					when "001010101111110" => rgb <= "101111";
					when "001010101111111" => rgb <= "101111";
					when "001010110000000" => rgb <= "101111";
					when "001010110000001" => rgb <= "101111";
					when "001010110000010" => rgb <= "101111";
					when "001010110000011" => rgb <= "101111";
					when "001010110000100" => rgb <= "101111";
					when "001010110000101" => rgb <= "101111";
					when "001010110000110" => rgb <= "101111";
					when "001010110000111" => rgb <= "101111";
					when "001010110001000" => rgb <= "101111";
					when "001010110001001" => rgb <= "101111";
					when "001010110001010" => rgb <= "101111";
					when "001010110001011" => rgb <= "101111";
					when "001010110001100" => rgb <= "101111";
					when "001010110001101" => rgb <= "101111";
					when "001010110001110" => rgb <= "101111";
					when "001010110001111" => rgb <= "101111";
					when "001010110010000" => rgb <= "101111";
					when "001010110010001" => rgb <= "101111";
					when "001010110010010" => rgb <= "101111";
					when "001010110010011" => rgb <= "101111";
					when "001010110010100" => rgb <= "101111";
					when "001010110010101" => rgb <= "101111";
					when "001010110010110" => rgb <= "101111";
					when "001010110010111" => rgb <= "101111";
					when "001010110011000" => rgb <= "101111";
					when "001010110011001" => rgb <= "101111";
					when "001010110011010" => rgb <= "101111";
					when "001010110011011" => rgb <= "101111";
					when "001010110011100" => rgb <= "101111";
					when "001010110011101" => rgb <= "101111";
					when "001010110011110" => rgb <= "101111";
					when "001010110011111" => rgb <= "101111";
					when "001011000000000" => rgb <= "001000";
					when "001011000000001" => rgb <= "001000";
					when "001011000000010" => rgb <= "001000";
					when "001011000000011" => rgb <= "001000";
					when "001011000000100" => rgb <= "001000";
					when "001011000000101" => rgb <= "001000";
					when "001011000000110" => rgb <= "001000";
					when "001011000000111" => rgb <= "001000";
					when "001011000001000" => rgb <= "001000";
					when "001011000001001" => rgb <= "001000";
					when "001011000001010" => rgb <= "001000";
					when "001011000001011" => rgb <= "001000";
					when "001011000001100" => rgb <= "001000";
					when "001011000001101" => rgb <= "001000";
					when "001011000001110" => rgb <= "001000";
					when "001011000001111" => rgb <= "001000";
					when "001011000010000" => rgb <= "001000";
					when "001011000010001" => rgb <= "001000";
					when "001011000010010" => rgb <= "001000";
					when "001011000010011" => rgb <= "001000";
					when "001011000010100" => rgb <= "001000";
					when "001011000010101" => rgb <= "001000";
					when "001011000010110" => rgb <= "001000";
					when "001011000010111" => rgb <= "001000";
					when "001011000011000" => rgb <= "001000";
					when "001011000011001" => rgb <= "001000";
					when "001011000011010" => rgb <= "001000";
					when "001011000011011" => rgb <= "001000";
					when "001011000011100" => rgb <= "001000";
					when "001011000011101" => rgb <= "001000";
					when "001011000011110" => rgb <= "001000";
					when "001011000011111" => rgb <= "001000";
					when "001011000100000" => rgb <= "001000";
					when "001011000100001" => rgb <= "001000";
					when "001011000100010" => rgb <= "001000";
					when "001011000100011" => rgb <= "001000";
					when "001011000100100" => rgb <= "001000";
					when "001011000100101" => rgb <= "001000";
					when "001011000100110" => rgb <= "001000";
					when "001011000100111" => rgb <= "001000";
					when "001011000101000" => rgb <= "001000";
					when "001011000101001" => rgb <= "001000";
					when "001011000101010" => rgb <= "001000";
					when "001011000101011" => rgb <= "001000";
					when "001011000101100" => rgb <= "001000";
					when "001011000101101" => rgb <= "001000";
					when "001011000101110" => rgb <= "001000";
					when "001011000101111" => rgb <= "001000";
					when "001011000110000" => rgb <= "001000";
					when "001011000110001" => rgb <= "001000";
					when "001011000110010" => rgb <= "001000";
					when "001011000110011" => rgb <= "001000";
					when "001011000110100" => rgb <= "001000";
					when "001011000110101" => rgb <= "001000";
					when "001011000110110" => rgb <= "001000";
					when "001011000110111" => rgb <= "001000";
					when "001011000111000" => rgb <= "001000";
					when "001011000111001" => rgb <= "001000";
					when "001011000111010" => rgb <= "001000";
					when "001011000111011" => rgb <= "001000";
					when "001011000111100" => rgb <= "001000";
					when "001011000111101" => rgb <= "001000";
					when "001011000111110" => rgb <= "001000";
					when "001011000111111" => rgb <= "001000";
					when "001011001000000" => rgb <= "001000";
					when "001011001000001" => rgb <= "001000";
					when "001011001000010" => rgb <= "001000";
					when "001011001000011" => rgb <= "001000";
					when "001011001000100" => rgb <= "001000";
					when "001011001000101" => rgb <= "001000";
					when "001011001000110" => rgb <= "001000";
					when "001011001000111" => rgb <= "001000";
					when "001011001001000" => rgb <= "001000";
					when "001011001001001" => rgb <= "001000";
					when "001011001001010" => rgb <= "001000";
					when "001011001001011" => rgb <= "001000";
					when "001011001001100" => rgb <= "001000";
					when "001011001001101" => rgb <= "001000";
					when "001011001001110" => rgb <= "001000";
					when "001011001001111" => rgb <= "001000";
					when "001011001010000" => rgb <= "000000";
					when "001011001010001" => rgb <= "000000";
					when "001011001010010" => rgb <= "000000";
					when "001011001010011" => rgb <= "000000";
					when "001011001010100" => rgb <= "101111";
					when "001011001010101" => rgb <= "101111";
					when "001011001010110" => rgb <= "101111";
					when "001011001010111" => rgb <= "101111";
					when "001011001011000" => rgb <= "101111";
					when "001011001011001" => rgb <= "101111";
					when "001011001011010" => rgb <= "101111";
					when "001011001011011" => rgb <= "101111";
					when "001011001011100" => rgb <= "101111";
					when "001011001011101" => rgb <= "101111";
					when "001011001011110" => rgb <= "101111";
					when "001011001011111" => rgb <= "101111";
					when "001011001100000" => rgb <= "101111";
					when "001011001100001" => rgb <= "101111";
					when "001011001100010" => rgb <= "101111";
					when "001011001100011" => rgb <= "101111";
					when "001011001100100" => rgb <= "101111";
					when "001011001100101" => rgb <= "101111";
					when "001011001100110" => rgb <= "101111";
					when "001011001100111" => rgb <= "101111";
					when "001011001101000" => rgb <= "101111";
					when "001011001101001" => rgb <= "101111";
					when "001011001101010" => rgb <= "101111";
					when "001011001101011" => rgb <= "101111";
					when "001011001101100" => rgb <= "101111";
					when "001011001101101" => rgb <= "101111";
					when "001011001101110" => rgb <= "101111";
					when "001011001101111" => rgb <= "101111";
					when "001011001110000" => rgb <= "101111";
					when "001011001110001" => rgb <= "101111";
					when "001011001110010" => rgb <= "101111";
					when "001011001110011" => rgb <= "101111";
					when "001011001110100" => rgb <= "101111";
					when "001011001110101" => rgb <= "101111";
					when "001011001110110" => rgb <= "101111";
					when "001011001110111" => rgb <= "101111";
					when "001011001111000" => rgb <= "101111";
					when "001011001111001" => rgb <= "101111";
					when "001011001111010" => rgb <= "101111";
					when "001011001111011" => rgb <= "101111";
					when "001011001111100" => rgb <= "101111";
					when "001011001111101" => rgb <= "101111";
					when "001011001111110" => rgb <= "101111";
					when "001011001111111" => rgb <= "101111";
					when "001011010000000" => rgb <= "101111";
					when "001011010000001" => rgb <= "101111";
					when "001011010000010" => rgb <= "101111";
					when "001011010000011" => rgb <= "101111";
					when "001011010000100" => rgb <= "101111";
					when "001011010000101" => rgb <= "101111";
					when "001011010000110" => rgb <= "101111";
					when "001011010000111" => rgb <= "101111";
					when "001011010001000" => rgb <= "101111";
					when "001011010001001" => rgb <= "101111";
					when "001011010001010" => rgb <= "101111";
					when "001011010001011" => rgb <= "101111";
					when "001011010001100" => rgb <= "101111";
					when "001011010001101" => rgb <= "101111";
					when "001011010001110" => rgb <= "101111";
					when "001011010001111" => rgb <= "101111";
					when "001011010010000" => rgb <= "101111";
					when "001011010010001" => rgb <= "101111";
					when "001011010010010" => rgb <= "101111";
					when "001011010010011" => rgb <= "101111";
					when "001011010010100" => rgb <= "101111";
					when "001011010010101" => rgb <= "101111";
					when "001011010010110" => rgb <= "101111";
					when "001011010010111" => rgb <= "101111";
					when "001011010011000" => rgb <= "101111";
					when "001011010011001" => rgb <= "101111";
					when "001011010011010" => rgb <= "101111";
					when "001011010011011" => rgb <= "101111";
					when "001011010011100" => rgb <= "101111";
					when "001011010011101" => rgb <= "101111";
					when "001011010011110" => rgb <= "101111";
					when "001011010011111" => rgb <= "101111";
					when "001011100000000" => rgb <= "001000";
					when "001011100000001" => rgb <= "001000";
					when "001011100000010" => rgb <= "001000";
					when "001011100000011" => rgb <= "001000";
					when "001011100000100" => rgb <= "001000";
					when "001011100000101" => rgb <= "001000";
					when "001011100000110" => rgb <= "001000";
					when "001011100000111" => rgb <= "001000";
					when "001011100001000" => rgb <= "001000";
					when "001011100001001" => rgb <= "001000";
					when "001011100001010" => rgb <= "001000";
					when "001011100001011" => rgb <= "001000";
					when "001011100001100" => rgb <= "001000";
					when "001011100001101" => rgb <= "001000";
					when "001011100001110" => rgb <= "001000";
					when "001011100001111" => rgb <= "001000";
					when "001011100010000" => rgb <= "001000";
					when "001011100010001" => rgb <= "001000";
					when "001011100010010" => rgb <= "001000";
					when "001011100010011" => rgb <= "001000";
					when "001011100010100" => rgb <= "001000";
					when "001011100010101" => rgb <= "001000";
					when "001011100010110" => rgb <= "001000";
					when "001011100010111" => rgb <= "001000";
					when "001011100011000" => rgb <= "001000";
					when "001011100011001" => rgb <= "001000";
					when "001011100011010" => rgb <= "001000";
					when "001011100011011" => rgb <= "001000";
					when "001011100011100" => rgb <= "001000";
					when "001011100011101" => rgb <= "001000";
					when "001011100011110" => rgb <= "001000";
					when "001011100011111" => rgb <= "001000";
					when "001011100100000" => rgb <= "001000";
					when "001011100100001" => rgb <= "001000";
					when "001011100100010" => rgb <= "001000";
					when "001011100100011" => rgb <= "001000";
					when "001011100100100" => rgb <= "001000";
					when "001011100100101" => rgb <= "001000";
					when "001011100100110" => rgb <= "001000";
					when "001011100100111" => rgb <= "001000";
					when "001011100101000" => rgb <= "001000";
					when "001011100101001" => rgb <= "001000";
					when "001011100101010" => rgb <= "001000";
					when "001011100101011" => rgb <= "001000";
					when "001011100101100" => rgb <= "001000";
					when "001011100101101" => rgb <= "001000";
					when "001011100101110" => rgb <= "001000";
					when "001011100101111" => rgb <= "001000";
					when "001011100110000" => rgb <= "001000";
					when "001011100110001" => rgb <= "001000";
					when "001011100110010" => rgb <= "001000";
					when "001011100110011" => rgb <= "001000";
					when "001011100110100" => rgb <= "001000";
					when "001011100110101" => rgb <= "001000";
					when "001011100110110" => rgb <= "001000";
					when "001011100110111" => rgb <= "001000";
					when "001011100111000" => rgb <= "001000";
					when "001011100111001" => rgb <= "001000";
					when "001011100111010" => rgb <= "001000";
					when "001011100111011" => rgb <= "001000";
					when "001011100111100" => rgb <= "001000";
					when "001011100111101" => rgb <= "001000";
					when "001011100111110" => rgb <= "001000";
					when "001011100111111" => rgb <= "001000";
					when "001011101000000" => rgb <= "001000";
					when "001011101000001" => rgb <= "001000";
					when "001011101000010" => rgb <= "001000";
					when "001011101000011" => rgb <= "001000";
					when "001011101000100" => rgb <= "001000";
					when "001011101000101" => rgb <= "001000";
					when "001011101000110" => rgb <= "001000";
					when "001011101000111" => rgb <= "001000";
					when "001011101001000" => rgb <= "001000";
					when "001011101001001" => rgb <= "001000";
					when "001011101001010" => rgb <= "001000";
					when "001011101001011" => rgb <= "001000";
					when "001011101001100" => rgb <= "001000";
					when "001011101001101" => rgb <= "001000";
					when "001011101001110" => rgb <= "001000";
					when "001011101001111" => rgb <= "001000";
					when "001011101010000" => rgb <= "000000";
					when "001011101010001" => rgb <= "000000";
					when "001011101010010" => rgb <= "000000";
					when "001011101010011" => rgb <= "000000";
					when "001011101010100" => rgb <= "101111";
					when "001011101010101" => rgb <= "101111";
					when "001011101010110" => rgb <= "101111";
					when "001011101010111" => rgb <= "101111";
					when "001011101011000" => rgb <= "101111";
					when "001011101011001" => rgb <= "101111";
					when "001011101011010" => rgb <= "101111";
					when "001011101011011" => rgb <= "101111";
					when "001011101011100" => rgb <= "101111";
					when "001011101011101" => rgb <= "101111";
					when "001011101011110" => rgb <= "101111";
					when "001011101011111" => rgb <= "101111";
					when "001011101100000" => rgb <= "101111";
					when "001011101100001" => rgb <= "101111";
					when "001011101100010" => rgb <= "101111";
					when "001011101100011" => rgb <= "101111";
					when "001011101100100" => rgb <= "101111";
					when "001011101100101" => rgb <= "101111";
					when "001011101100110" => rgb <= "101111";
					when "001011101100111" => rgb <= "101111";
					when "001011101101000" => rgb <= "101111";
					when "001011101101001" => rgb <= "101111";
					when "001011101101010" => rgb <= "101111";
					when "001011101101011" => rgb <= "101111";
					when "001011101101100" => rgb <= "101111";
					when "001011101101101" => rgb <= "101111";
					when "001011101101110" => rgb <= "101111";
					when "001011101101111" => rgb <= "101111";
					when "001011101110000" => rgb <= "101111";
					when "001011101110001" => rgb <= "101111";
					when "001011101110010" => rgb <= "101111";
					when "001011101110011" => rgb <= "101111";
					when "001011101110100" => rgb <= "101111";
					when "001011101110101" => rgb <= "101111";
					when "001011101110110" => rgb <= "101111";
					when "001011101110111" => rgb <= "101111";
					when "001011101111000" => rgb <= "101111";
					when "001011101111001" => rgb <= "101111";
					when "001011101111010" => rgb <= "101111";
					when "001011101111011" => rgb <= "101111";
					when "001011101111100" => rgb <= "101111";
					when "001011101111101" => rgb <= "101111";
					when "001011101111110" => rgb <= "101111";
					when "001011101111111" => rgb <= "101111";
					when "001011110000000" => rgb <= "101111";
					when "001011110000001" => rgb <= "101111";
					when "001011110000010" => rgb <= "101111";
					when "001011110000011" => rgb <= "101111";
					when "001011110000100" => rgb <= "101111";
					when "001011110000101" => rgb <= "101111";
					when "001011110000110" => rgb <= "101111";
					when "001011110000111" => rgb <= "101111";
					when "001011110001000" => rgb <= "101111";
					when "001011110001001" => rgb <= "101111";
					when "001011110001010" => rgb <= "101111";
					when "001011110001011" => rgb <= "101111";
					when "001011110001100" => rgb <= "101111";
					when "001011110001101" => rgb <= "101111";
					when "001011110001110" => rgb <= "101111";
					when "001011110001111" => rgb <= "101111";
					when "001011110010000" => rgb <= "101111";
					when "001011110010001" => rgb <= "101111";
					when "001011110010010" => rgb <= "101111";
					when "001011110010011" => rgb <= "101111";
					when "001011110010100" => rgb <= "101111";
					when "001011110010101" => rgb <= "101111";
					when "001011110010110" => rgb <= "101111";
					when "001011110010111" => rgb <= "101111";
					when "001011110011000" => rgb <= "101111";
					when "001011110011001" => rgb <= "101111";
					when "001011110011010" => rgb <= "101111";
					when "001011110011011" => rgb <= "101111";
					when "001011110011100" => rgb <= "101111";
					when "001011110011101" => rgb <= "101111";
					when "001011110011110" => rgb <= "101111";
					when "001011110011111" => rgb <= "101111";
					when "001100000000000" => rgb <= "001000";
					when "001100000000001" => rgb <= "001000";
					when "001100000000010" => rgb <= "001000";
					when "001100000000011" => rgb <= "001000";
					when "001100000000100" => rgb <= "001000";
					when "001100000000101" => rgb <= "001000";
					when "001100000000110" => rgb <= "001000";
					when "001100000000111" => rgb <= "001000";
					when "001100000001000" => rgb <= "001000";
					when "001100000001001" => rgb <= "001000";
					when "001100000001010" => rgb <= "001000";
					when "001100000001011" => rgb <= "001000";
					when "001100000001100" => rgb <= "001000";
					when "001100000001101" => rgb <= "001000";
					when "001100000001110" => rgb <= "001000";
					when "001100000001111" => rgb <= "001000";
					when "001100000010000" => rgb <= "001000";
					when "001100000010001" => rgb <= "001000";
					when "001100000010010" => rgb <= "001000";
					when "001100000010011" => rgb <= "001000";
					when "001100000010100" => rgb <= "001000";
					when "001100000010101" => rgb <= "001000";
					when "001100000010110" => rgb <= "001000";
					when "001100000010111" => rgb <= "001000";
					when "001100000011000" => rgb <= "001000";
					when "001100000011001" => rgb <= "001000";
					when "001100000011010" => rgb <= "001000";
					when "001100000011011" => rgb <= "001000";
					when "001100000011100" => rgb <= "001000";
					when "001100000011101" => rgb <= "001000";
					when "001100000011110" => rgb <= "001000";
					when "001100000011111" => rgb <= "001000";
					when "001100000100000" => rgb <= "001000";
					when "001100000100001" => rgb <= "001000";
					when "001100000100010" => rgb <= "001000";
					when "001100000100011" => rgb <= "001000";
					when "001100000100100" => rgb <= "001000";
					when "001100000100101" => rgb <= "001000";
					when "001100000100110" => rgb <= "001000";
					when "001100000100111" => rgb <= "001000";
					when "001100000101000" => rgb <= "001000";
					when "001100000101001" => rgb <= "001000";
					when "001100000101010" => rgb <= "001000";
					when "001100000101011" => rgb <= "001000";
					when "001100000101100" => rgb <= "001000";
					when "001100000101101" => rgb <= "001000";
					when "001100000101110" => rgb <= "001000";
					when "001100000101111" => rgb <= "001000";
					when "001100000110000" => rgb <= "001000";
					when "001100000110001" => rgb <= "001000";
					when "001100000110010" => rgb <= "001000";
					when "001100000110011" => rgb <= "001000";
					when "001100000110100" => rgb <= "001000";
					when "001100000110101" => rgb <= "001000";
					when "001100000110110" => rgb <= "001000";
					when "001100000110111" => rgb <= "001000";
					when "001100000111000" => rgb <= "001000";
					when "001100000111001" => rgb <= "001000";
					when "001100000111010" => rgb <= "001000";
					when "001100000111011" => rgb <= "001000";
					when "001100000111100" => rgb <= "001000";
					when "001100000111101" => rgb <= "001000";
					when "001100000111110" => rgb <= "001000";
					when "001100000111111" => rgb <= "001000";
					when "001100001000000" => rgb <= "001000";
					when "001100001000001" => rgb <= "001000";
					when "001100001000010" => rgb <= "001000";
					when "001100001000011" => rgb <= "001000";
					when "001100001000100" => rgb <= "001000";
					when "001100001000101" => rgb <= "001000";
					when "001100001000110" => rgb <= "001000";
					when "001100001000111" => rgb <= "001000";
					when "001100001001000" => rgb <= "001000";
					when "001100001001001" => rgb <= "001000";
					when "001100001001010" => rgb <= "001000";
					when "001100001001011" => rgb <= "001000";
					when "001100001001100" => rgb <= "001000";
					when "001100001001101" => rgb <= "001000";
					when "001100001001110" => rgb <= "001000";
					when "001100001001111" => rgb <= "001000";
					when "001100001010000" => rgb <= "001000";
					when "001100001010001" => rgb <= "001000";
					when "001100001010010" => rgb <= "000000";
					when "001100001010011" => rgb <= "000000";
					when "001100001010100" => rgb <= "000000";
					when "001100001010101" => rgb <= "000000";
					when "001100001010110" => rgb <= "101111";
					when "001100001010111" => rgb <= "101111";
					when "001100001011000" => rgb <= "101111";
					when "001100001011001" => rgb <= "101111";
					when "001100001011010" => rgb <= "101111";
					when "001100001011011" => rgb <= "101111";
					when "001100001011100" => rgb <= "101111";
					when "001100001011101" => rgb <= "101111";
					when "001100001011110" => rgb <= "101111";
					when "001100001011111" => rgb <= "101111";
					when "001100001100000" => rgb <= "101111";
					when "001100001100001" => rgb <= "101111";
					when "001100001100010" => rgb <= "101111";
					when "001100001100011" => rgb <= "101111";
					when "001100001100100" => rgb <= "101111";
					when "001100001100101" => rgb <= "101111";
					when "001100001100110" => rgb <= "101111";
					when "001100001100111" => rgb <= "101111";
					when "001100001101000" => rgb <= "101111";
					when "001100001101001" => rgb <= "101111";
					when "001100001101010" => rgb <= "101111";
					when "001100001101011" => rgb <= "101111";
					when "001100001101100" => rgb <= "101111";
					when "001100001101101" => rgb <= "101111";
					when "001100001101110" => rgb <= "101111";
					when "001100001101111" => rgb <= "101111";
					when "001100001110000" => rgb <= "101111";
					when "001100001110001" => rgb <= "101111";
					when "001100001110010" => rgb <= "101111";
					when "001100001110011" => rgb <= "101111";
					when "001100001110100" => rgb <= "101111";
					when "001100001110101" => rgb <= "101111";
					when "001100001110110" => rgb <= "101111";
					when "001100001110111" => rgb <= "101111";
					when "001100001111000" => rgb <= "101111";
					when "001100001111001" => rgb <= "101111";
					when "001100001111010" => rgb <= "101111";
					when "001100001111011" => rgb <= "101111";
					when "001100001111100" => rgb <= "101111";
					when "001100001111101" => rgb <= "101111";
					when "001100001111110" => rgb <= "101111";
					when "001100001111111" => rgb <= "101111";
					when "001100010000000" => rgb <= "101111";
					when "001100010000001" => rgb <= "101111";
					when "001100010000010" => rgb <= "101111";
					when "001100010000011" => rgb <= "101111";
					when "001100010000100" => rgb <= "101111";
					when "001100010000101" => rgb <= "101111";
					when "001100010000110" => rgb <= "101111";
					when "001100010000111" => rgb <= "101111";
					when "001100010001000" => rgb <= "101111";
					when "001100010001001" => rgb <= "101111";
					when "001100010001010" => rgb <= "101111";
					when "001100010001011" => rgb <= "101111";
					when "001100010001100" => rgb <= "101111";
					when "001100010001101" => rgb <= "101111";
					when "001100010001110" => rgb <= "101111";
					when "001100010001111" => rgb <= "101111";
					when "001100010010000" => rgb <= "101111";
					when "001100010010001" => rgb <= "101111";
					when "001100010010010" => rgb <= "101111";
					when "001100010010011" => rgb <= "101111";
					when "001100010010100" => rgb <= "101111";
					when "001100010010101" => rgb <= "101111";
					when "001100010010110" => rgb <= "101111";
					when "001100010010111" => rgb <= "101111";
					when "001100010011000" => rgb <= "101111";
					when "001100010011001" => rgb <= "101111";
					when "001100010011010" => rgb <= "101111";
					when "001100010011011" => rgb <= "101111";
					when "001100010011100" => rgb <= "101111";
					when "001100010011101" => rgb <= "101111";
					when "001100010011110" => rgb <= "101111";
					when "001100010011111" => rgb <= "101111";
					when "001100100000000" => rgb <= "001000";
					when "001100100000001" => rgb <= "001000";
					when "001100100000010" => rgb <= "001000";
					when "001100100000011" => rgb <= "001000";
					when "001100100000100" => rgb <= "001000";
					when "001100100000101" => rgb <= "001000";
					when "001100100000110" => rgb <= "001000";
					when "001100100000111" => rgb <= "001000";
					when "001100100001000" => rgb <= "001000";
					when "001100100001001" => rgb <= "001000";
					when "001100100001010" => rgb <= "001000";
					when "001100100001011" => rgb <= "001000";
					when "001100100001100" => rgb <= "001000";
					when "001100100001101" => rgb <= "001000";
					when "001100100001110" => rgb <= "001000";
					when "001100100001111" => rgb <= "001000";
					when "001100100010000" => rgb <= "001000";
					when "001100100010001" => rgb <= "001000";
					when "001100100010010" => rgb <= "001000";
					when "001100100010011" => rgb <= "001000";
					when "001100100010100" => rgb <= "001000";
					when "001100100010101" => rgb <= "001000";
					when "001100100010110" => rgb <= "001000";
					when "001100100010111" => rgb <= "001000";
					when "001100100011000" => rgb <= "001000";
					when "001100100011001" => rgb <= "001000";
					when "001100100011010" => rgb <= "001000";
					when "001100100011011" => rgb <= "001000";
					when "001100100011100" => rgb <= "001000";
					when "001100100011101" => rgb <= "001000";
					when "001100100011110" => rgb <= "001000";
					when "001100100011111" => rgb <= "001000";
					when "001100100100000" => rgb <= "001000";
					when "001100100100001" => rgb <= "001000";
					when "001100100100010" => rgb <= "001000";
					when "001100100100011" => rgb <= "001000";
					when "001100100100100" => rgb <= "001000";
					when "001100100100101" => rgb <= "001000";
					when "001100100100110" => rgb <= "001000";
					when "001100100100111" => rgb <= "001000";
					when "001100100101000" => rgb <= "001000";
					when "001100100101001" => rgb <= "001000";
					when "001100100101010" => rgb <= "001000";
					when "001100100101011" => rgb <= "001000";
					when "001100100101100" => rgb <= "001000";
					when "001100100101101" => rgb <= "001000";
					when "001100100101110" => rgb <= "001000";
					when "001100100101111" => rgb <= "001000";
					when "001100100110000" => rgb <= "001000";
					when "001100100110001" => rgb <= "001000";
					when "001100100110010" => rgb <= "001000";
					when "001100100110011" => rgb <= "001000";
					when "001100100110100" => rgb <= "001000";
					when "001100100110101" => rgb <= "001000";
					when "001100100110110" => rgb <= "001000";
					when "001100100110111" => rgb <= "001000";
					when "001100100111000" => rgb <= "001000";
					when "001100100111001" => rgb <= "001000";
					when "001100100111010" => rgb <= "001000";
					when "001100100111011" => rgb <= "001000";
					when "001100100111100" => rgb <= "001000";
					when "001100100111101" => rgb <= "001000";
					when "001100100111110" => rgb <= "001000";
					when "001100100111111" => rgb <= "001000";
					when "001100101000000" => rgb <= "001000";
					when "001100101000001" => rgb <= "001000";
					when "001100101000010" => rgb <= "001000";
					when "001100101000011" => rgb <= "001000";
					when "001100101000100" => rgb <= "001000";
					when "001100101000101" => rgb <= "001000";
					when "001100101000110" => rgb <= "001000";
					when "001100101000111" => rgb <= "001000";
					when "001100101001000" => rgb <= "001000";
					when "001100101001001" => rgb <= "001000";
					when "001100101001010" => rgb <= "001000";
					when "001100101001011" => rgb <= "001000";
					when "001100101001100" => rgb <= "001000";
					when "001100101001101" => rgb <= "001000";
					when "001100101001110" => rgb <= "001000";
					when "001100101001111" => rgb <= "001000";
					when "001100101010000" => rgb <= "001000";
					when "001100101010001" => rgb <= "001000";
					when "001100101010010" => rgb <= "000000";
					when "001100101010011" => rgb <= "000000";
					when "001100101010100" => rgb <= "000000";
					when "001100101010101" => rgb <= "000000";
					when "001100101010110" => rgb <= "101111";
					when "001100101010111" => rgb <= "101111";
					when "001100101011000" => rgb <= "101111";
					when "001100101011001" => rgb <= "101111";
					when "001100101011010" => rgb <= "101111";
					when "001100101011011" => rgb <= "101111";
					when "001100101011100" => rgb <= "101111";
					when "001100101011101" => rgb <= "101111";
					when "001100101011110" => rgb <= "101111";
					when "001100101011111" => rgb <= "101111";
					when "001100101100000" => rgb <= "101111";
					when "001100101100001" => rgb <= "101111";
					when "001100101100010" => rgb <= "101111";
					when "001100101100011" => rgb <= "101111";
					when "001100101100100" => rgb <= "101111";
					when "001100101100101" => rgb <= "101111";
					when "001100101100110" => rgb <= "101111";
					when "001100101100111" => rgb <= "101111";
					when "001100101101000" => rgb <= "101111";
					when "001100101101001" => rgb <= "101111";
					when "001100101101010" => rgb <= "101111";
					when "001100101101011" => rgb <= "101111";
					when "001100101101100" => rgb <= "101111";
					when "001100101101101" => rgb <= "101111";
					when "001100101101110" => rgb <= "101111";
					when "001100101101111" => rgb <= "101111";
					when "001100101110000" => rgb <= "101111";
					when "001100101110001" => rgb <= "101111";
					when "001100101110010" => rgb <= "101111";
					when "001100101110011" => rgb <= "101111";
					when "001100101110100" => rgb <= "101111";
					when "001100101110101" => rgb <= "101111";
					when "001100101110110" => rgb <= "101111";
					when "001100101110111" => rgb <= "101111";
					when "001100101111000" => rgb <= "101111";
					when "001100101111001" => rgb <= "101111";
					when "001100101111010" => rgb <= "101111";
					when "001100101111011" => rgb <= "101111";
					when "001100101111100" => rgb <= "101111";
					when "001100101111101" => rgb <= "101111";
					when "001100101111110" => rgb <= "101111";
					when "001100101111111" => rgb <= "101111";
					when "001100110000000" => rgb <= "101111";
					when "001100110000001" => rgb <= "101111";
					when "001100110000010" => rgb <= "101111";
					when "001100110000011" => rgb <= "101111";
					when "001100110000100" => rgb <= "101111";
					when "001100110000101" => rgb <= "101111";
					when "001100110000110" => rgb <= "101111";
					when "001100110000111" => rgb <= "101111";
					when "001100110001000" => rgb <= "101111";
					when "001100110001001" => rgb <= "101111";
					when "001100110001010" => rgb <= "101111";
					when "001100110001011" => rgb <= "101111";
					when "001100110001100" => rgb <= "101111";
					when "001100110001101" => rgb <= "101111";
					when "001100110001110" => rgb <= "101111";
					when "001100110001111" => rgb <= "101111";
					when "001100110010000" => rgb <= "101111";
					when "001100110010001" => rgb <= "101111";
					when "001100110010010" => rgb <= "101111";
					when "001100110010011" => rgb <= "101111";
					when "001100110010100" => rgb <= "101111";
					when "001100110010101" => rgb <= "101111";
					when "001100110010110" => rgb <= "101111";
					when "001100110010111" => rgb <= "101111";
					when "001100110011000" => rgb <= "101111";
					when "001100110011001" => rgb <= "101111";
					when "001100110011010" => rgb <= "101111";
					when "001100110011011" => rgb <= "101111";
					when "001100110011100" => rgb <= "101111";
					when "001100110011101" => rgb <= "101111";
					when "001100110011110" => rgb <= "101111";
					when "001100110011111" => rgb <= "101111";
					when "001101000000000" => rgb <= "001000";
					when "001101000000001" => rgb <= "001000";
					when "001101000000010" => rgb <= "001000";
					when "001101000000011" => rgb <= "001000";
					when "001101000000100" => rgb <= "001000";
					when "001101000000101" => rgb <= "001000";
					when "001101000000110" => rgb <= "001000";
					when "001101000000111" => rgb <= "001000";
					when "001101000001000" => rgb <= "001000";
					when "001101000001001" => rgb <= "001000";
					when "001101000001010" => rgb <= "001000";
					when "001101000001011" => rgb <= "001000";
					when "001101000001100" => rgb <= "001000";
					when "001101000001101" => rgb <= "001000";
					when "001101000001110" => rgb <= "001000";
					when "001101000001111" => rgb <= "001000";
					when "001101000010000" => rgb <= "001000";
					when "001101000010001" => rgb <= "001000";
					when "001101000010010" => rgb <= "001000";
					when "001101000010011" => rgb <= "001000";
					when "001101000010100" => rgb <= "001000";
					when "001101000010101" => rgb <= "001000";
					when "001101000010110" => rgb <= "001000";
					when "001101000010111" => rgb <= "001000";
					when "001101000011000" => rgb <= "001000";
					when "001101000011001" => rgb <= "001000";
					when "001101000011010" => rgb <= "001000";
					when "001101000011011" => rgb <= "001000";
					when "001101000011100" => rgb <= "001000";
					when "001101000011101" => rgb <= "001000";
					when "001101000011110" => rgb <= "001000";
					when "001101000011111" => rgb <= "001000";
					when "001101000100000" => rgb <= "001000";
					when "001101000100001" => rgb <= "001000";
					when "001101000100010" => rgb <= "001000";
					when "001101000100011" => rgb <= "001000";
					when "001101000100100" => rgb <= "001000";
					when "001101000100101" => rgb <= "001000";
					when "001101000100110" => rgb <= "001000";
					when "001101000100111" => rgb <= "001000";
					when "001101000101000" => rgb <= "001000";
					when "001101000101001" => rgb <= "001000";
					when "001101000101010" => rgb <= "001000";
					when "001101000101011" => rgb <= "001000";
					when "001101000101100" => rgb <= "001000";
					when "001101000101101" => rgb <= "001000";
					when "001101000101110" => rgb <= "001000";
					when "001101000101111" => rgb <= "001000";
					when "001101000110000" => rgb <= "001000";
					when "001101000110001" => rgb <= "001000";
					when "001101000110010" => rgb <= "001000";
					when "001101000110011" => rgb <= "001000";
					when "001101000110100" => rgb <= "001000";
					when "001101000110101" => rgb <= "001000";
					when "001101000110110" => rgb <= "001000";
					when "001101000110111" => rgb <= "001000";
					when "001101000111000" => rgb <= "001000";
					when "001101000111001" => rgb <= "001000";
					when "001101000111010" => rgb <= "001000";
					when "001101000111011" => rgb <= "001000";
					when "001101000111100" => rgb <= "001000";
					when "001101000111101" => rgb <= "001000";
					when "001101000111110" => rgb <= "001000";
					when "001101000111111" => rgb <= "001000";
					when "001101001000000" => rgb <= "001000";
					when "001101001000001" => rgb <= "001000";
					when "001101001000010" => rgb <= "001000";
					when "001101001000011" => rgb <= "001000";
					when "001101001000100" => rgb <= "001000";
					when "001101001000101" => rgb <= "001000";
					when "001101001000110" => rgb <= "001000";
					when "001101001000111" => rgb <= "001000";
					when "001101001001000" => rgb <= "001000";
					when "001101001001001" => rgb <= "001000";
					when "001101001001010" => rgb <= "001000";
					when "001101001001011" => rgb <= "001000";
					when "001101001001100" => rgb <= "001000";
					when "001101001001101" => rgb <= "001000";
					when "001101001001110" => rgb <= "001000";
					when "001101001001111" => rgb <= "001000";
					when "001101001010000" => rgb <= "001000";
					when "001101001010001" => rgb <= "001000";
					when "001101001010010" => rgb <= "001000";
					when "001101001010011" => rgb <= "001000";
					when "001101001010100" => rgb <= "000000";
					when "001101001010101" => rgb <= "000000";
					when "001101001010110" => rgb <= "101111";
					when "001101001010111" => rgb <= "101111";
					when "001101001011000" => rgb <= "101111";
					when "001101001011001" => rgb <= "101111";
					when "001101001011010" => rgb <= "101111";
					when "001101001011011" => rgb <= "101111";
					when "001101001011100" => rgb <= "101111";
					when "001101001011101" => rgb <= "101111";
					when "001101001011110" => rgb <= "101111";
					when "001101001011111" => rgb <= "101111";
					when "001101001100000" => rgb <= "101111";
					when "001101001100001" => rgb <= "101111";
					when "001101001100010" => rgb <= "101111";
					when "001101001100011" => rgb <= "101111";
					when "001101001100100" => rgb <= "101111";
					when "001101001100101" => rgb <= "101111";
					when "001101001100110" => rgb <= "101111";
					when "001101001100111" => rgb <= "101111";
					when "001101001101000" => rgb <= "101111";
					when "001101001101001" => rgb <= "101111";
					when "001101001101010" => rgb <= "101111";
					when "001101001101011" => rgb <= "101111";
					when "001101001101100" => rgb <= "101111";
					when "001101001101101" => rgb <= "101111";
					when "001101001101110" => rgb <= "101111";
					when "001101001101111" => rgb <= "101111";
					when "001101001110000" => rgb <= "101111";
					when "001101001110001" => rgb <= "101111";
					when "001101001110010" => rgb <= "101111";
					when "001101001110011" => rgb <= "101111";
					when "001101001110100" => rgb <= "101111";
					when "001101001110101" => rgb <= "101111";
					when "001101001110110" => rgb <= "101111";
					when "001101001110111" => rgb <= "101111";
					when "001101001111000" => rgb <= "101111";
					when "001101001111001" => rgb <= "101111";
					when "001101001111010" => rgb <= "101111";
					when "001101001111011" => rgb <= "101111";
					when "001101001111100" => rgb <= "101111";
					when "001101001111101" => rgb <= "101111";
					when "001101001111110" => rgb <= "101111";
					when "001101001111111" => rgb <= "101111";
					when "001101010000000" => rgb <= "101111";
					when "001101010000001" => rgb <= "101111";
					when "001101010000010" => rgb <= "101111";
					when "001101010000011" => rgb <= "101111";
					when "001101010000100" => rgb <= "101111";
					when "001101010000101" => rgb <= "101111";
					when "001101010000110" => rgb <= "101111";
					when "001101010000111" => rgb <= "101111";
					when "001101010001000" => rgb <= "101111";
					when "001101010001001" => rgb <= "101111";
					when "001101010001010" => rgb <= "101111";
					when "001101010001011" => rgb <= "101111";
					when "001101010001100" => rgb <= "101111";
					when "001101010001101" => rgb <= "101111";
					when "001101010001110" => rgb <= "101111";
					when "001101010001111" => rgb <= "101111";
					when "001101010010000" => rgb <= "101111";
					when "001101010010001" => rgb <= "101111";
					when "001101010010010" => rgb <= "101111";
					when "001101010010011" => rgb <= "101111";
					when "001101010010100" => rgb <= "101111";
					when "001101010010101" => rgb <= "101111";
					when "001101010010110" => rgb <= "101111";
					when "001101010010111" => rgb <= "101111";
					when "001101010011000" => rgb <= "101111";
					when "001101010011001" => rgb <= "101111";
					when "001101010011010" => rgb <= "101111";
					when "001101010011011" => rgb <= "101111";
					when "001101010011100" => rgb <= "101111";
					when "001101010011101" => rgb <= "101111";
					when "001101010011110" => rgb <= "101111";
					when "001101010011111" => rgb <= "101111";
					when "001101100000000" => rgb <= "001000";
					when "001101100000001" => rgb <= "001000";
					when "001101100000010" => rgb <= "001000";
					when "001101100000011" => rgb <= "001000";
					when "001101100000100" => rgb <= "001000";
					when "001101100000101" => rgb <= "001000";
					when "001101100000110" => rgb <= "001000";
					when "001101100000111" => rgb <= "001000";
					when "001101100001000" => rgb <= "001000";
					when "001101100001001" => rgb <= "001000";
					when "001101100001010" => rgb <= "001000";
					when "001101100001011" => rgb <= "001000";
					when "001101100001100" => rgb <= "001000";
					when "001101100001101" => rgb <= "001000";
					when "001101100001110" => rgb <= "001000";
					when "001101100001111" => rgb <= "001000";
					when "001101100010000" => rgb <= "001000";
					when "001101100010001" => rgb <= "001000";
					when "001101100010010" => rgb <= "001000";
					when "001101100010011" => rgb <= "001000";
					when "001101100010100" => rgb <= "001000";
					when "001101100010101" => rgb <= "001000";
					when "001101100010110" => rgb <= "001000";
					when "001101100010111" => rgb <= "001000";
					when "001101100011000" => rgb <= "001000";
					when "001101100011001" => rgb <= "001000";
					when "001101100011010" => rgb <= "001000";
					when "001101100011011" => rgb <= "001000";
					when "001101100011100" => rgb <= "001000";
					when "001101100011101" => rgb <= "001000";
					when "001101100011110" => rgb <= "001000";
					when "001101100011111" => rgb <= "001000";
					when "001101100100000" => rgb <= "001000";
					when "001101100100001" => rgb <= "001000";
					when "001101100100010" => rgb <= "001000";
					when "001101100100011" => rgb <= "001000";
					when "001101100100100" => rgb <= "001000";
					when "001101100100101" => rgb <= "001000";
					when "001101100100110" => rgb <= "001000";
					when "001101100100111" => rgb <= "001000";
					when "001101100101000" => rgb <= "001000";
					when "001101100101001" => rgb <= "001000";
					when "001101100101010" => rgb <= "001000";
					when "001101100101011" => rgb <= "001000";
					when "001101100101100" => rgb <= "001000";
					when "001101100101101" => rgb <= "001000";
					when "001101100101110" => rgb <= "001000";
					when "001101100101111" => rgb <= "001000";
					when "001101100110000" => rgb <= "001000";
					when "001101100110001" => rgb <= "001000";
					when "001101100110010" => rgb <= "001000";
					when "001101100110011" => rgb <= "001000";
					when "001101100110100" => rgb <= "001000";
					when "001101100110101" => rgb <= "001000";
					when "001101100110110" => rgb <= "001000";
					when "001101100110111" => rgb <= "001000";
					when "001101100111000" => rgb <= "001000";
					when "001101100111001" => rgb <= "001000";
					when "001101100111010" => rgb <= "001000";
					when "001101100111011" => rgb <= "001000";
					when "001101100111100" => rgb <= "001000";
					when "001101100111101" => rgb <= "001000";
					when "001101100111110" => rgb <= "001000";
					when "001101100111111" => rgb <= "001000";
					when "001101101000000" => rgb <= "001000";
					when "001101101000001" => rgb <= "001000";
					when "001101101000010" => rgb <= "001000";
					when "001101101000011" => rgb <= "001000";
					when "001101101000100" => rgb <= "001000";
					when "001101101000101" => rgb <= "001000";
					when "001101101000110" => rgb <= "001000";
					when "001101101000111" => rgb <= "001000";
					when "001101101001000" => rgb <= "001000";
					when "001101101001001" => rgb <= "001000";
					when "001101101001010" => rgb <= "001000";
					when "001101101001011" => rgb <= "001000";
					when "001101101001100" => rgb <= "001000";
					when "001101101001101" => rgb <= "001000";
					when "001101101001110" => rgb <= "001000";
					when "001101101001111" => rgb <= "001000";
					when "001101101010000" => rgb <= "001000";
					when "001101101010001" => rgb <= "001000";
					when "001101101010010" => rgb <= "001000";
					when "001101101010011" => rgb <= "001000";
					when "001101101010100" => rgb <= "000000";
					when "001101101010101" => rgb <= "000000";
					when "001101101010110" => rgb <= "101111";
					when "001101101010111" => rgb <= "101111";
					when "001101101011000" => rgb <= "101111";
					when "001101101011001" => rgb <= "101111";
					when "001101101011010" => rgb <= "101111";
					when "001101101011011" => rgb <= "101111";
					when "001101101011100" => rgb <= "101111";
					when "001101101011101" => rgb <= "101111";
					when "001101101011110" => rgb <= "101111";
					when "001101101011111" => rgb <= "101111";
					when "001101101100000" => rgb <= "101111";
					when "001101101100001" => rgb <= "101111";
					when "001101101100010" => rgb <= "101111";
					when "001101101100011" => rgb <= "101111";
					when "001101101100100" => rgb <= "101111";
					when "001101101100101" => rgb <= "101111";
					when "001101101100110" => rgb <= "101111";
					when "001101101100111" => rgb <= "101111";
					when "001101101101000" => rgb <= "101111";
					when "001101101101001" => rgb <= "101111";
					when "001101101101010" => rgb <= "101111";
					when "001101101101011" => rgb <= "101111";
					when "001101101101100" => rgb <= "101111";
					when "001101101101101" => rgb <= "101111";
					when "001101101101110" => rgb <= "101111";
					when "001101101101111" => rgb <= "101111";
					when "001101101110000" => rgb <= "101111";
					when "001101101110001" => rgb <= "101111";
					when "001101101110010" => rgb <= "101111";
					when "001101101110011" => rgb <= "101111";
					when "001101101110100" => rgb <= "101111";
					when "001101101110101" => rgb <= "101111";
					when "001101101110110" => rgb <= "101111";
					when "001101101110111" => rgb <= "101111";
					when "001101101111000" => rgb <= "101111";
					when "001101101111001" => rgb <= "101111";
					when "001101101111010" => rgb <= "101111";
					when "001101101111011" => rgb <= "101111";
					when "001101101111100" => rgb <= "101111";
					when "001101101111101" => rgb <= "101111";
					when "001101101111110" => rgb <= "101111";
					when "001101101111111" => rgb <= "101111";
					when "001101110000000" => rgb <= "101111";
					when "001101110000001" => rgb <= "101111";
					when "001101110000010" => rgb <= "101111";
					when "001101110000011" => rgb <= "101111";
					when "001101110000100" => rgb <= "101111";
					when "001101110000101" => rgb <= "101111";
					when "001101110000110" => rgb <= "101111";
					when "001101110000111" => rgb <= "101111";
					when "001101110001000" => rgb <= "101111";
					when "001101110001001" => rgb <= "101111";
					when "001101110001010" => rgb <= "101111";
					when "001101110001011" => rgb <= "101111";
					when "001101110001100" => rgb <= "101111";
					when "001101110001101" => rgb <= "101111";
					when "001101110001110" => rgb <= "101111";
					when "001101110001111" => rgb <= "101111";
					when "001101110010000" => rgb <= "101111";
					when "001101110010001" => rgb <= "101111";
					when "001101110010010" => rgb <= "101111";
					when "001101110010011" => rgb <= "101111";
					when "001101110010100" => rgb <= "101111";
					when "001101110010101" => rgb <= "101111";
					when "001101110010110" => rgb <= "101111";
					when "001101110010111" => rgb <= "101111";
					when "001101110011000" => rgb <= "101111";
					when "001101110011001" => rgb <= "101111";
					when "001101110011010" => rgb <= "101111";
					when "001101110011011" => rgb <= "101111";
					when "001101110011100" => rgb <= "101111";
					when "001101110011101" => rgb <= "101111";
					when "001101110011110" => rgb <= "101111";
					when "001101110011111" => rgb <= "101111";
					when "001110000000000" => rgb <= "001000";
					when "001110000000001" => rgb <= "001000";
					when "001110000000010" => rgb <= "001000";
					when "001110000000011" => rgb <= "001000";
					when "001110000000100" => rgb <= "001000";
					when "001110000000101" => rgb <= "001000";
					when "001110000000110" => rgb <= "001000";
					when "001110000000111" => rgb <= "001000";
					when "001110000001000" => rgb <= "001000";
					when "001110000001001" => rgb <= "001000";
					when "001110000001010" => rgb <= "001000";
					when "001110000001011" => rgb <= "001000";
					when "001110000001100" => rgb <= "001000";
					when "001110000001101" => rgb <= "001000";
					when "001110000001110" => rgb <= "001000";
					when "001110000001111" => rgb <= "001000";
					when "001110000010000" => rgb <= "001000";
					when "001110000010001" => rgb <= "001000";
					when "001110000010010" => rgb <= "001000";
					when "001110000010011" => rgb <= "001000";
					when "001110000010100" => rgb <= "001000";
					when "001110000010101" => rgb <= "001000";
					when "001110000010110" => rgb <= "001000";
					when "001110000010111" => rgb <= "001000";
					when "001110000011000" => rgb <= "001000";
					when "001110000011001" => rgb <= "001000";
					when "001110000011010" => rgb <= "001000";
					when "001110000011011" => rgb <= "001000";
					when "001110000011100" => rgb <= "001000";
					when "001110000011101" => rgb <= "001000";
					when "001110000011110" => rgb <= "001000";
					when "001110000011111" => rgb <= "001000";
					when "001110000100000" => rgb <= "001000";
					when "001110000100001" => rgb <= "001000";
					when "001110000100010" => rgb <= "001000";
					when "001110000100011" => rgb <= "001000";
					when "001110000100100" => rgb <= "001000";
					when "001110000100101" => rgb <= "001000";
					when "001110000100110" => rgb <= "001000";
					when "001110000100111" => rgb <= "001000";
					when "001110000101000" => rgb <= "001000";
					when "001110000101001" => rgb <= "001000";
					when "001110000101010" => rgb <= "001000";
					when "001110000101011" => rgb <= "001000";
					when "001110000101100" => rgb <= "001000";
					when "001110000101101" => rgb <= "001000";
					when "001110000101110" => rgb <= "001000";
					when "001110000101111" => rgb <= "001000";
					when "001110000110000" => rgb <= "001000";
					when "001110000110001" => rgb <= "001000";
					when "001110000110010" => rgb <= "001000";
					when "001110000110011" => rgb <= "001000";
					when "001110000110100" => rgb <= "001000";
					when "001110000110101" => rgb <= "001000";
					when "001110000110110" => rgb <= "001000";
					when "001110000110111" => rgb <= "001000";
					when "001110000111000" => rgb <= "001000";
					when "001110000111001" => rgb <= "001000";
					when "001110000111010" => rgb <= "001000";
					when "001110000111011" => rgb <= "001000";
					when "001110000111100" => rgb <= "001000";
					when "001110000111101" => rgb <= "001000";
					when "001110000111110" => rgb <= "001000";
					when "001110000111111" => rgb <= "001000";
					when "001110001000000" => rgb <= "001000";
					when "001110001000001" => rgb <= "001000";
					when "001110001000010" => rgb <= "001000";
					when "001110001000011" => rgb <= "001000";
					when "001110001000100" => rgb <= "001000";
					when "001110001000101" => rgb <= "001000";
					when "001110001000110" => rgb <= "001000";
					when "001110001000111" => rgb <= "001000";
					when "001110001001000" => rgb <= "001000";
					when "001110001001001" => rgb <= "001000";
					when "001110001001010" => rgb <= "001000";
					when "001110001001011" => rgb <= "001000";
					when "001110001001100" => rgb <= "001000";
					when "001110001001101" => rgb <= "001000";
					when "001110001001110" => rgb <= "001000";
					when "001110001001111" => rgb <= "001000";
					when "001110001010000" => rgb <= "001000";
					when "001110001010001" => rgb <= "001000";
					when "001110001010010" => rgb <= "001000";
					when "001110001010011" => rgb <= "001000";
					when "001110001010100" => rgb <= "000000";
					when "001110001010101" => rgb <= "000000";
					when "001110001010110" => rgb <= "000000";
					when "001110001010111" => rgb <= "000000";
					when "001110001011000" => rgb <= "101111";
					when "001110001011001" => rgb <= "101111";
					when "001110001011010" => rgb <= "101111";
					when "001110001011011" => rgb <= "101111";
					when "001110001011100" => rgb <= "101111";
					when "001110001011101" => rgb <= "101111";
					when "001110001011110" => rgb <= "101111";
					when "001110001011111" => rgb <= "101111";
					when "001110001100000" => rgb <= "101111";
					when "001110001100001" => rgb <= "101111";
					when "001110001100010" => rgb <= "101111";
					when "001110001100011" => rgb <= "101111";
					when "001110001100100" => rgb <= "101111";
					when "001110001100101" => rgb <= "101111";
					when "001110001100110" => rgb <= "101111";
					when "001110001100111" => rgb <= "101111";
					when "001110001101000" => rgb <= "101111";
					when "001110001101001" => rgb <= "101111";
					when "001110001101010" => rgb <= "101111";
					when "001110001101011" => rgb <= "101111";
					when "001110001101100" => rgb <= "101111";
					when "001110001101101" => rgb <= "101111";
					when "001110001101110" => rgb <= "101111";
					when "001110001101111" => rgb <= "101111";
					when "001110001110000" => rgb <= "101111";
					when "001110001110001" => rgb <= "101111";
					when "001110001110010" => rgb <= "101111";
					when "001110001110011" => rgb <= "101111";
					when "001110001110100" => rgb <= "101111";
					when "001110001110101" => rgb <= "101111";
					when "001110001110110" => rgb <= "101111";
					when "001110001110111" => rgb <= "101111";
					when "001110001111000" => rgb <= "101111";
					when "001110001111001" => rgb <= "101111";
					when "001110001111010" => rgb <= "101111";
					when "001110001111011" => rgb <= "101111";
					when "001110001111100" => rgb <= "101111";
					when "001110001111101" => rgb <= "101111";
					when "001110001111110" => rgb <= "101111";
					when "001110001111111" => rgb <= "101111";
					when "001110010000000" => rgb <= "101111";
					when "001110010000001" => rgb <= "101111";
					when "001110010000010" => rgb <= "101111";
					when "001110010000011" => rgb <= "101111";
					when "001110010000100" => rgb <= "101111";
					when "001110010000101" => rgb <= "101111";
					when "001110010000110" => rgb <= "101111";
					when "001110010000111" => rgb <= "101111";
					when "001110010001000" => rgb <= "101111";
					when "001110010001001" => rgb <= "101111";
					when "001110010001010" => rgb <= "101111";
					when "001110010001011" => rgb <= "101111";
					when "001110010001100" => rgb <= "101111";
					when "001110010001101" => rgb <= "101111";
					when "001110010001110" => rgb <= "101111";
					when "001110010001111" => rgb <= "101111";
					when "001110010010000" => rgb <= "101111";
					when "001110010010001" => rgb <= "101111";
					when "001110010010010" => rgb <= "101111";
					when "001110010010011" => rgb <= "101111";
					when "001110010010100" => rgb <= "101111";
					when "001110010010101" => rgb <= "101111";
					when "001110010010110" => rgb <= "101111";
					when "001110010010111" => rgb <= "101111";
					when "001110010011000" => rgb <= "101111";
					when "001110010011001" => rgb <= "101111";
					when "001110010011010" => rgb <= "101111";
					when "001110010011011" => rgb <= "101111";
					when "001110010011100" => rgb <= "101111";
					when "001110010011101" => rgb <= "101111";
					when "001110010011110" => rgb <= "101111";
					when "001110010011111" => rgb <= "101111";
					when "001110100000000" => rgb <= "001000";
					when "001110100000001" => rgb <= "001000";
					when "001110100000010" => rgb <= "001000";
					when "001110100000011" => rgb <= "001000";
					when "001110100000100" => rgb <= "001000";
					when "001110100000101" => rgb <= "001000";
					when "001110100000110" => rgb <= "001000";
					when "001110100000111" => rgb <= "001000";
					when "001110100001000" => rgb <= "001000";
					when "001110100001001" => rgb <= "001000";
					when "001110100001010" => rgb <= "001000";
					when "001110100001011" => rgb <= "001000";
					when "001110100001100" => rgb <= "001000";
					when "001110100001101" => rgb <= "001000";
					when "001110100001110" => rgb <= "001000";
					when "001110100001111" => rgb <= "001000";
					when "001110100010000" => rgb <= "001000";
					when "001110100010001" => rgb <= "001000";
					when "001110100010010" => rgb <= "001000";
					when "001110100010011" => rgb <= "001000";
					when "001110100010100" => rgb <= "001000";
					when "001110100010101" => rgb <= "001000";
					when "001110100010110" => rgb <= "001000";
					when "001110100010111" => rgb <= "001000";
					when "001110100011000" => rgb <= "001000";
					when "001110100011001" => rgb <= "001000";
					when "001110100011010" => rgb <= "001000";
					when "001110100011011" => rgb <= "001000";
					when "001110100011100" => rgb <= "001000";
					when "001110100011101" => rgb <= "001000";
					when "001110100011110" => rgb <= "001000";
					when "001110100011111" => rgb <= "001000";
					when "001110100100000" => rgb <= "001000";
					when "001110100100001" => rgb <= "001000";
					when "001110100100010" => rgb <= "001000";
					when "001110100100011" => rgb <= "001000";
					when "001110100100100" => rgb <= "001000";
					when "001110100100101" => rgb <= "001000";
					when "001110100100110" => rgb <= "001000";
					when "001110100100111" => rgb <= "001000";
					when "001110100101000" => rgb <= "001000";
					when "001110100101001" => rgb <= "001000";
					when "001110100101010" => rgb <= "001000";
					when "001110100101011" => rgb <= "001000";
					when "001110100101100" => rgb <= "001000";
					when "001110100101101" => rgb <= "001000";
					when "001110100101110" => rgb <= "001000";
					when "001110100101111" => rgb <= "001000";
					when "001110100110000" => rgb <= "001000";
					when "001110100110001" => rgb <= "001000";
					when "001110100110010" => rgb <= "001000";
					when "001110100110011" => rgb <= "001000";
					when "001110100110100" => rgb <= "001000";
					when "001110100110101" => rgb <= "001000";
					when "001110100110110" => rgb <= "001000";
					when "001110100110111" => rgb <= "001000";
					when "001110100111000" => rgb <= "001000";
					when "001110100111001" => rgb <= "001000";
					when "001110100111010" => rgb <= "001000";
					when "001110100111011" => rgb <= "001000";
					when "001110100111100" => rgb <= "001000";
					when "001110100111101" => rgb <= "001000";
					when "001110100111110" => rgb <= "001000";
					when "001110100111111" => rgb <= "001000";
					when "001110101000000" => rgb <= "001000";
					when "001110101000001" => rgb <= "001000";
					when "001110101000010" => rgb <= "001000";
					when "001110101000011" => rgb <= "001000";
					when "001110101000100" => rgb <= "001000";
					when "001110101000101" => rgb <= "001000";
					when "001110101000110" => rgb <= "001000";
					when "001110101000111" => rgb <= "001000";
					when "001110101001000" => rgb <= "001000";
					when "001110101001001" => rgb <= "001000";
					when "001110101001010" => rgb <= "001000";
					when "001110101001011" => rgb <= "001000";
					when "001110101001100" => rgb <= "001000";
					when "001110101001101" => rgb <= "001000";
					when "001110101001110" => rgb <= "001000";
					when "001110101001111" => rgb <= "001000";
					when "001110101010000" => rgb <= "001000";
					when "001110101010001" => rgb <= "001000";
					when "001110101010010" => rgb <= "001000";
					when "001110101010011" => rgb <= "001000";
					when "001110101010100" => rgb <= "000000";
					when "001110101010101" => rgb <= "000000";
					when "001110101010110" => rgb <= "000000";
					when "001110101010111" => rgb <= "000000";
					when "001110101011000" => rgb <= "101111";
					when "001110101011001" => rgb <= "101111";
					when "001110101011010" => rgb <= "101111";
					when "001110101011011" => rgb <= "101111";
					when "001110101011100" => rgb <= "101111";
					when "001110101011101" => rgb <= "101111";
					when "001110101011110" => rgb <= "101111";
					when "001110101011111" => rgb <= "101111";
					when "001110101100000" => rgb <= "101111";
					when "001110101100001" => rgb <= "101111";
					when "001110101100010" => rgb <= "101111";
					when "001110101100011" => rgb <= "101111";
					when "001110101100100" => rgb <= "101111";
					when "001110101100101" => rgb <= "101111";
					when "001110101100110" => rgb <= "101111";
					when "001110101100111" => rgb <= "101111";
					when "001110101101000" => rgb <= "101111";
					when "001110101101001" => rgb <= "101111";
					when "001110101101010" => rgb <= "101111";
					when "001110101101011" => rgb <= "101111";
					when "001110101101100" => rgb <= "101111";
					when "001110101101101" => rgb <= "101111";
					when "001110101101110" => rgb <= "101111";
					when "001110101101111" => rgb <= "101111";
					when "001110101110000" => rgb <= "101111";
					when "001110101110001" => rgb <= "101111";
					when "001110101110010" => rgb <= "101111";
					when "001110101110011" => rgb <= "101111";
					when "001110101110100" => rgb <= "101111";
					when "001110101110101" => rgb <= "101111";
					when "001110101110110" => rgb <= "101111";
					when "001110101110111" => rgb <= "101111";
					when "001110101111000" => rgb <= "101111";
					when "001110101111001" => rgb <= "101111";
					when "001110101111010" => rgb <= "101111";
					when "001110101111011" => rgb <= "101111";
					when "001110101111100" => rgb <= "101111";
					when "001110101111101" => rgb <= "101111";
					when "001110101111110" => rgb <= "101111";
					when "001110101111111" => rgb <= "101111";
					when "001110110000000" => rgb <= "101111";
					when "001110110000001" => rgb <= "101111";
					when "001110110000010" => rgb <= "101111";
					when "001110110000011" => rgb <= "101111";
					when "001110110000100" => rgb <= "101111";
					when "001110110000101" => rgb <= "101111";
					when "001110110000110" => rgb <= "101111";
					when "001110110000111" => rgb <= "101111";
					when "001110110001000" => rgb <= "101111";
					when "001110110001001" => rgb <= "101111";
					when "001110110001010" => rgb <= "101111";
					when "001110110001011" => rgb <= "101111";
					when "001110110001100" => rgb <= "101111";
					when "001110110001101" => rgb <= "101111";
					when "001110110001110" => rgb <= "101111";
					when "001110110001111" => rgb <= "101111";
					when "001110110010000" => rgb <= "101111";
					when "001110110010001" => rgb <= "101111";
					when "001110110010010" => rgb <= "101111";
					when "001110110010011" => rgb <= "101111";
					when "001110110010100" => rgb <= "101111";
					when "001110110010101" => rgb <= "101111";
					when "001110110010110" => rgb <= "101111";
					when "001110110010111" => rgb <= "101111";
					when "001110110011000" => rgb <= "101111";
					when "001110110011001" => rgb <= "101111";
					when "001110110011010" => rgb <= "101111";
					when "001110110011011" => rgb <= "101111";
					when "001110110011100" => rgb <= "101111";
					when "001110110011101" => rgb <= "101111";
					when "001110110011110" => rgb <= "101111";
					when "001110110011111" => rgb <= "101111";
					when "001111000000000" => rgb <= "001000";
					when "001111000000001" => rgb <= "001000";
					when "001111000000010" => rgb <= "001000";
					when "001111000000011" => rgb <= "001000";
					when "001111000000100" => rgb <= "001000";
					when "001111000000101" => rgb <= "001000";
					when "001111000000110" => rgb <= "001000";
					when "001111000000111" => rgb <= "001000";
					when "001111000001000" => rgb <= "001000";
					when "001111000001001" => rgb <= "001000";
					when "001111000001010" => rgb <= "001000";
					when "001111000001011" => rgb <= "001000";
					when "001111000001100" => rgb <= "001000";
					when "001111000001101" => rgb <= "001000";
					when "001111000001110" => rgb <= "001000";
					when "001111000001111" => rgb <= "001000";
					when "001111000010000" => rgb <= "001000";
					when "001111000010001" => rgb <= "001000";
					when "001111000010010" => rgb <= "001000";
					when "001111000010011" => rgb <= "001000";
					when "001111000010100" => rgb <= "001000";
					when "001111000010101" => rgb <= "001000";
					when "001111000010110" => rgb <= "001000";
					when "001111000010111" => rgb <= "001000";
					when "001111000011000" => rgb <= "001000";
					when "001111000011001" => rgb <= "001000";
					when "001111000011010" => rgb <= "001000";
					when "001111000011011" => rgb <= "001000";
					when "001111000011100" => rgb <= "001000";
					when "001111000011101" => rgb <= "001000";
					when "001111000011110" => rgb <= "001000";
					when "001111000011111" => rgb <= "001000";
					when "001111000100000" => rgb <= "001000";
					when "001111000100001" => rgb <= "001000";
					when "001111000100010" => rgb <= "001000";
					when "001111000100011" => rgb <= "001000";
					when "001111000100100" => rgb <= "001000";
					when "001111000100101" => rgb <= "001000";
					when "001111000100110" => rgb <= "001000";
					when "001111000100111" => rgb <= "001000";
					when "001111000101000" => rgb <= "001000";
					when "001111000101001" => rgb <= "001000";
					when "001111000101010" => rgb <= "001000";
					when "001111000101011" => rgb <= "001000";
					when "001111000101100" => rgb <= "001000";
					when "001111000101101" => rgb <= "001000";
					when "001111000101110" => rgb <= "001000";
					when "001111000101111" => rgb <= "001000";
					when "001111000110000" => rgb <= "001000";
					when "001111000110001" => rgb <= "001000";
					when "001111000110010" => rgb <= "001000";
					when "001111000110011" => rgb <= "001000";
					when "001111000110100" => rgb <= "001000";
					when "001111000110101" => rgb <= "001000";
					when "001111000110110" => rgb <= "001000";
					when "001111000110111" => rgb <= "001000";
					when "001111000111000" => rgb <= "001000";
					when "001111000111001" => rgb <= "001000";
					when "001111000111010" => rgb <= "001000";
					when "001111000111011" => rgb <= "001000";
					when "001111000111100" => rgb <= "001000";
					when "001111000111101" => rgb <= "001000";
					when "001111000111110" => rgb <= "001000";
					when "001111000111111" => rgb <= "001000";
					when "001111001000000" => rgb <= "001000";
					when "001111001000001" => rgb <= "001000";
					when "001111001000010" => rgb <= "001000";
					when "001111001000011" => rgb <= "001000";
					when "001111001000100" => rgb <= "001000";
					when "001111001000101" => rgb <= "001000";
					when "001111001000110" => rgb <= "001000";
					when "001111001000111" => rgb <= "001000";
					when "001111001001000" => rgb <= "001000";
					when "001111001001001" => rgb <= "001000";
					when "001111001001010" => rgb <= "001000";
					when "001111001001011" => rgb <= "001000";
					when "001111001001100" => rgb <= "001000";
					when "001111001001101" => rgb <= "001000";
					when "001111001001110" => rgb <= "001000";
					when "001111001001111" => rgb <= "001000";
					when "001111001010000" => rgb <= "001000";
					when "001111001010001" => rgb <= "001000";
					when "001111001010010" => rgb <= "001000";
					when "001111001010011" => rgb <= "001000";
					when "001111001010100" => rgb <= "001000";
					when "001111001010101" => rgb <= "001000";
					when "001111001010110" => rgb <= "000000";
					when "001111001010111" => rgb <= "000000";
					when "001111001011000" => rgb <= "000000";
					when "001111001011001" => rgb <= "000000";
					when "001111001011010" => rgb <= "101111";
					when "001111001011011" => rgb <= "101111";
					when "001111001011100" => rgb <= "101111";
					when "001111001011101" => rgb <= "101111";
					when "001111001011110" => rgb <= "101111";
					when "001111001011111" => rgb <= "101111";
					when "001111001100000" => rgb <= "101111";
					when "001111001100001" => rgb <= "101111";
					when "001111001100010" => rgb <= "101111";
					when "001111001100011" => rgb <= "101111";
					when "001111001100100" => rgb <= "101111";
					when "001111001100101" => rgb <= "101111";
					when "001111001100110" => rgb <= "101111";
					when "001111001100111" => rgb <= "101111";
					when "001111001101000" => rgb <= "101111";
					when "001111001101001" => rgb <= "101111";
					when "001111001101010" => rgb <= "101111";
					when "001111001101011" => rgb <= "101111";
					when "001111001101100" => rgb <= "101111";
					when "001111001101101" => rgb <= "101111";
					when "001111001101110" => rgb <= "101111";
					when "001111001101111" => rgb <= "101111";
					when "001111001110000" => rgb <= "101111";
					when "001111001110001" => rgb <= "101111";
					when "001111001110010" => rgb <= "101111";
					when "001111001110011" => rgb <= "101111";
					when "001111001110100" => rgb <= "101111";
					when "001111001110101" => rgb <= "101111";
					when "001111001110110" => rgb <= "101111";
					when "001111001110111" => rgb <= "101111";
					when "001111001111000" => rgb <= "101111";
					when "001111001111001" => rgb <= "101111";
					when "001111001111010" => rgb <= "101111";
					when "001111001111011" => rgb <= "101111";
					when "001111001111100" => rgb <= "101111";
					when "001111001111101" => rgb <= "101111";
					when "001111001111110" => rgb <= "101111";
					when "001111001111111" => rgb <= "101111";
					when "001111010000000" => rgb <= "101111";
					when "001111010000001" => rgb <= "101111";
					when "001111010000010" => rgb <= "101111";
					when "001111010000011" => rgb <= "101111";
					when "001111010000100" => rgb <= "101111";
					when "001111010000101" => rgb <= "101111";
					when "001111010000110" => rgb <= "101111";
					when "001111010000111" => rgb <= "101111";
					when "001111010001000" => rgb <= "101111";
					when "001111010001001" => rgb <= "101111";
					when "001111010001010" => rgb <= "101111";
					when "001111010001011" => rgb <= "101111";
					when "001111010001100" => rgb <= "101111";
					when "001111010001101" => rgb <= "101111";
					when "001111010001110" => rgb <= "101111";
					when "001111010001111" => rgb <= "101111";
					when "001111010010000" => rgb <= "101111";
					when "001111010010001" => rgb <= "101111";
					when "001111010010010" => rgb <= "101111";
					when "001111010010011" => rgb <= "101111";
					when "001111010010100" => rgb <= "101111";
					when "001111010010101" => rgb <= "101111";
					when "001111010010110" => rgb <= "101111";
					when "001111010010111" => rgb <= "101111";
					when "001111010011000" => rgb <= "101111";
					when "001111010011001" => rgb <= "101111";
					when "001111010011010" => rgb <= "101111";
					when "001111010011011" => rgb <= "101111";
					when "001111010011100" => rgb <= "101111";
					when "001111010011101" => rgb <= "101111";
					when "001111010011110" => rgb <= "101111";
					when "001111010011111" => rgb <= "101111";
					when "001111100000000" => rgb <= "001000";
					when "001111100000001" => rgb <= "001000";
					when "001111100000010" => rgb <= "001000";
					when "001111100000011" => rgb <= "001000";
					when "001111100000100" => rgb <= "001000";
					when "001111100000101" => rgb <= "001000";
					when "001111100000110" => rgb <= "001000";
					when "001111100000111" => rgb <= "001000";
					when "001111100001000" => rgb <= "001000";
					when "001111100001001" => rgb <= "001000";
					when "001111100001010" => rgb <= "001000";
					when "001111100001011" => rgb <= "001000";
					when "001111100001100" => rgb <= "001000";
					when "001111100001101" => rgb <= "001000";
					when "001111100001110" => rgb <= "001000";
					when "001111100001111" => rgb <= "001000";
					when "001111100010000" => rgb <= "001000";
					when "001111100010001" => rgb <= "001000";
					when "001111100010010" => rgb <= "001000";
					when "001111100010011" => rgb <= "001000";
					when "001111100010100" => rgb <= "001000";
					when "001111100010101" => rgb <= "001000";
					when "001111100010110" => rgb <= "001000";
					when "001111100010111" => rgb <= "001000";
					when "001111100011000" => rgb <= "001000";
					when "001111100011001" => rgb <= "001000";
					when "001111100011010" => rgb <= "001000";
					when "001111100011011" => rgb <= "001000";
					when "001111100011100" => rgb <= "001000";
					when "001111100011101" => rgb <= "001000";
					when "001111100011110" => rgb <= "001000";
					when "001111100011111" => rgb <= "001000";
					when "001111100100000" => rgb <= "001000";
					when "001111100100001" => rgb <= "001000";
					when "001111100100010" => rgb <= "001000";
					when "001111100100011" => rgb <= "001000";
					when "001111100100100" => rgb <= "001000";
					when "001111100100101" => rgb <= "001000";
					when "001111100100110" => rgb <= "001000";
					when "001111100100111" => rgb <= "001000";
					when "001111100101000" => rgb <= "001000";
					when "001111100101001" => rgb <= "001000";
					when "001111100101010" => rgb <= "001000";
					when "001111100101011" => rgb <= "001000";
					when "001111100101100" => rgb <= "001000";
					when "001111100101101" => rgb <= "001000";
					when "001111100101110" => rgb <= "001000";
					when "001111100101111" => rgb <= "001000";
					when "001111100110000" => rgb <= "001000";
					when "001111100110001" => rgb <= "001000";
					when "001111100110010" => rgb <= "001000";
					when "001111100110011" => rgb <= "001000";
					when "001111100110100" => rgb <= "001000";
					when "001111100110101" => rgb <= "001000";
					when "001111100110110" => rgb <= "001000";
					when "001111100110111" => rgb <= "001000";
					when "001111100111000" => rgb <= "001000";
					when "001111100111001" => rgb <= "001000";
					when "001111100111010" => rgb <= "001000";
					when "001111100111011" => rgb <= "001000";
					when "001111100111100" => rgb <= "001000";
					when "001111100111101" => rgb <= "001000";
					when "001111100111110" => rgb <= "001000";
					when "001111100111111" => rgb <= "001000";
					when "001111101000000" => rgb <= "001000";
					when "001111101000001" => rgb <= "001000";
					when "001111101000010" => rgb <= "001000";
					when "001111101000011" => rgb <= "001000";
					when "001111101000100" => rgb <= "001000";
					when "001111101000101" => rgb <= "001000";
					when "001111101000110" => rgb <= "001000";
					when "001111101000111" => rgb <= "001000";
					when "001111101001000" => rgb <= "001000";
					when "001111101001001" => rgb <= "001000";
					when "001111101001010" => rgb <= "001000";
					when "001111101001011" => rgb <= "001000";
					when "001111101001100" => rgb <= "001000";
					when "001111101001101" => rgb <= "001000";
					when "001111101001110" => rgb <= "001000";
					when "001111101001111" => rgb <= "001000";
					when "001111101010000" => rgb <= "001000";
					when "001111101010001" => rgb <= "001000";
					when "001111101010010" => rgb <= "001000";
					when "001111101010011" => rgb <= "001000";
					when "001111101010100" => rgb <= "001000";
					when "001111101010101" => rgb <= "001000";
					when "001111101010110" => rgb <= "000000";
					when "001111101010111" => rgb <= "000000";
					when "001111101011000" => rgb <= "000000";
					when "001111101011001" => rgb <= "000000";
					when "001111101011010" => rgb <= "101111";
					when "001111101011011" => rgb <= "101111";
					when "001111101011100" => rgb <= "101111";
					when "001111101011101" => rgb <= "101111";
					when "001111101011110" => rgb <= "101111";
					when "001111101011111" => rgb <= "101111";
					when "001111101100000" => rgb <= "101111";
					when "001111101100001" => rgb <= "101111";
					when "001111101100010" => rgb <= "101111";
					when "001111101100011" => rgb <= "101111";
					when "001111101100100" => rgb <= "101111";
					when "001111101100101" => rgb <= "101111";
					when "001111101100110" => rgb <= "101111";
					when "001111101100111" => rgb <= "101111";
					when "001111101101000" => rgb <= "101111";
					when "001111101101001" => rgb <= "101111";
					when "001111101101010" => rgb <= "101111";
					when "001111101101011" => rgb <= "101111";
					when "001111101101100" => rgb <= "101111";
					when "001111101101101" => rgb <= "101111";
					when "001111101101110" => rgb <= "101111";
					when "001111101101111" => rgb <= "101111";
					when "001111101110000" => rgb <= "101111";
					when "001111101110001" => rgb <= "101111";
					when "001111101110010" => rgb <= "101111";
					when "001111101110011" => rgb <= "101111";
					when "001111101110100" => rgb <= "101111";
					when "001111101110101" => rgb <= "101111";
					when "001111101110110" => rgb <= "101111";
					when "001111101110111" => rgb <= "101111";
					when "001111101111000" => rgb <= "101111";
					when "001111101111001" => rgb <= "101111";
					when "001111101111010" => rgb <= "101111";
					when "001111101111011" => rgb <= "101111";
					when "001111101111100" => rgb <= "101111";
					when "001111101111101" => rgb <= "101111";
					when "001111101111110" => rgb <= "101111";
					when "001111101111111" => rgb <= "101111";
					when "001111110000000" => rgb <= "101111";
					when "001111110000001" => rgb <= "101111";
					when "001111110000010" => rgb <= "101111";
					when "001111110000011" => rgb <= "101111";
					when "001111110000100" => rgb <= "101111";
					when "001111110000101" => rgb <= "101111";
					when "001111110000110" => rgb <= "101111";
					when "001111110000111" => rgb <= "101111";
					when "001111110001000" => rgb <= "101111";
					when "001111110001001" => rgb <= "101111";
					when "001111110001010" => rgb <= "101111";
					when "001111110001011" => rgb <= "101111";
					when "001111110001100" => rgb <= "101111";
					when "001111110001101" => rgb <= "101111";
					when "001111110001110" => rgb <= "101111";
					when "001111110001111" => rgb <= "101111";
					when "001111110010000" => rgb <= "101111";
					when "001111110010001" => rgb <= "101111";
					when "001111110010010" => rgb <= "101111";
					when "001111110010011" => rgb <= "101111";
					when "001111110010100" => rgb <= "101111";
					when "001111110010101" => rgb <= "101111";
					when "001111110010110" => rgb <= "101111";
					when "001111110010111" => rgb <= "101111";
					when "001111110011000" => rgb <= "101111";
					when "001111110011001" => rgb <= "101111";
					when "001111110011010" => rgb <= "101111";
					when "001111110011011" => rgb <= "101111";
					when "001111110011100" => rgb <= "101111";
					when "001111110011101" => rgb <= "101111";
					when "001111110011110" => rgb <= "101111";
					when "001111110011111" => rgb <= "101111";
					when "010000000000000" => rgb <= "001000";
					when "010000000000001" => rgb <= "001000";
					when "010000000000010" => rgb <= "001000";
					when "010000000000011" => rgb <= "001000";
					when "010000000000100" => rgb <= "001000";
					when "010000000000101" => rgb <= "001000";
					when "010000000000110" => rgb <= "001000";
					when "010000000000111" => rgb <= "001000";
					when "010000000001000" => rgb <= "001000";
					when "010000000001001" => rgb <= "001000";
					when "010000000001010" => rgb <= "001000";
					when "010000000001011" => rgb <= "001000";
					when "010000000001100" => rgb <= "001000";
					when "010000000001101" => rgb <= "001000";
					when "010000000001110" => rgb <= "001000";
					when "010000000001111" => rgb <= "001000";
					when "010000000010000" => rgb <= "001000";
					when "010000000010001" => rgb <= "001000";
					when "010000000010010" => rgb <= "001000";
					when "010000000010011" => rgb <= "001000";
					when "010000000010100" => rgb <= "001000";
					when "010000000010101" => rgb <= "001000";
					when "010000000010110" => rgb <= "001000";
					when "010000000010111" => rgb <= "001000";
					when "010000000011000" => rgb <= "001000";
					when "010000000011001" => rgb <= "001000";
					when "010000000011010" => rgb <= "001000";
					when "010000000011011" => rgb <= "001000";
					when "010000000011100" => rgb <= "001000";
					when "010000000011101" => rgb <= "001000";
					when "010000000011110" => rgb <= "001000";
					when "010000000011111" => rgb <= "001000";
					when "010000000100000" => rgb <= "001000";
					when "010000000100001" => rgb <= "001000";
					when "010000000100010" => rgb <= "001000";
					when "010000000100011" => rgb <= "001000";
					when "010000000100100" => rgb <= "001000";
					when "010000000100101" => rgb <= "001000";
					when "010000000100110" => rgb <= "001000";
					when "010000000100111" => rgb <= "001000";
					when "010000000101000" => rgb <= "001000";
					when "010000000101001" => rgb <= "001000";
					when "010000000101010" => rgb <= "001000";
					when "010000000101011" => rgb <= "001000";
					when "010000000101100" => rgb <= "001000";
					when "010000000101101" => rgb <= "001000";
					when "010000000101110" => rgb <= "001000";
					when "010000000101111" => rgb <= "001000";
					when "010000000110000" => rgb <= "001000";
					when "010000000110001" => rgb <= "001000";
					when "010000000110010" => rgb <= "001000";
					when "010000000110011" => rgb <= "001000";
					when "010000000110100" => rgb <= "001000";
					when "010000000110101" => rgb <= "001000";
					when "010000000110110" => rgb <= "001000";
					when "010000000110111" => rgb <= "001000";
					when "010000000111000" => rgb <= "001000";
					when "010000000111001" => rgb <= "001000";
					when "010000000111010" => rgb <= "001000";
					when "010000000111011" => rgb <= "001000";
					when "010000000111100" => rgb <= "001000";
					when "010000000111101" => rgb <= "001000";
					when "010000000111110" => rgb <= "001000";
					when "010000000111111" => rgb <= "001000";
					when "010000001000000" => rgb <= "001000";
					when "010000001000001" => rgb <= "001000";
					when "010000001000010" => rgb <= "001000";
					when "010000001000011" => rgb <= "001000";
					when "010000001000100" => rgb <= "001000";
					when "010000001000101" => rgb <= "001000";
					when "010000001000110" => rgb <= "001000";
					when "010000001000111" => rgb <= "001000";
					when "010000001001000" => rgb <= "001000";
					when "010000001001001" => rgb <= "001000";
					when "010000001001010" => rgb <= "001000";
					when "010000001001011" => rgb <= "001000";
					when "010000001001100" => rgb <= "001000";
					when "010000001001101" => rgb <= "001000";
					when "010000001001110" => rgb <= "001000";
					when "010000001001111" => rgb <= "001000";
					when "010000001010000" => rgb <= "001000";
					when "010000001010001" => rgb <= "001000";
					when "010000001010010" => rgb <= "001000";
					when "010000001010011" => rgb <= "001000";
					when "010000001010100" => rgb <= "001000";
					when "010000001010101" => rgb <= "001000";
					when "010000001010110" => rgb <= "001000";
					when "010000001010111" => rgb <= "001000";
					when "010000001011000" => rgb <= "001000";
					when "010000001011001" => rgb <= "001000";
					when "010000001011010" => rgb <= "000000";
					when "010000001011011" => rgb <= "000000";
					when "010000001011100" => rgb <= "101111";
					when "010000001011101" => rgb <= "101111";
					when "010000001011110" => rgb <= "101111";
					when "010000001011111" => rgb <= "101111";
					when "010000001100000" => rgb <= "101111";
					when "010000001100001" => rgb <= "101111";
					when "010000001100010" => rgb <= "101111";
					when "010000001100011" => rgb <= "101111";
					when "010000001100100" => rgb <= "101111";
					when "010000001100101" => rgb <= "101111";
					when "010000001100110" => rgb <= "101111";
					when "010000001100111" => rgb <= "101111";
					when "010000001101000" => rgb <= "101111";
					when "010000001101001" => rgb <= "101111";
					when "010000001101010" => rgb <= "101111";
					when "010000001101011" => rgb <= "101111";
					when "010000001101100" => rgb <= "101111";
					when "010000001101101" => rgb <= "101111";
					when "010000001101110" => rgb <= "101111";
					when "010000001101111" => rgb <= "101111";
					when "010000001110000" => rgb <= "101111";
					when "010000001110001" => rgb <= "101111";
					when "010000001110010" => rgb <= "101111";
					when "010000001110011" => rgb <= "101111";
					when "010000001110100" => rgb <= "101111";
					when "010000001110101" => rgb <= "101111";
					when "010000001110110" => rgb <= "101111";
					when "010000001110111" => rgb <= "101111";
					when "010000001111000" => rgb <= "101111";
					when "010000001111001" => rgb <= "101111";
					when "010000001111010" => rgb <= "101111";
					when "010000001111011" => rgb <= "101111";
					when "010000001111100" => rgb <= "101111";
					when "010000001111101" => rgb <= "101111";
					when "010000001111110" => rgb <= "101111";
					when "010000001111111" => rgb <= "101111";
					when "010000010000000" => rgb <= "101111";
					when "010000010000001" => rgb <= "101111";
					when "010000010000010" => rgb <= "101111";
					when "010000010000011" => rgb <= "101111";
					when "010000010000100" => rgb <= "101111";
					when "010000010000101" => rgb <= "101111";
					when "010000010000110" => rgb <= "101111";
					when "010000010000111" => rgb <= "101111";
					when "010000010001000" => rgb <= "101111";
					when "010000010001001" => rgb <= "101111";
					when "010000010001010" => rgb <= "101111";
					when "010000010001011" => rgb <= "101111";
					when "010000010001100" => rgb <= "101111";
					when "010000010001101" => rgb <= "101111";
					when "010000010001110" => rgb <= "101111";
					when "010000010001111" => rgb <= "101111";
					when "010000010010000" => rgb <= "101111";
					when "010000010010001" => rgb <= "101111";
					when "010000010010010" => rgb <= "101111";
					when "010000010010011" => rgb <= "101111";
					when "010000010010100" => rgb <= "101111";
					when "010000010010101" => rgb <= "101111";
					when "010000010010110" => rgb <= "101111";
					when "010000010010111" => rgb <= "101111";
					when "010000010011000" => rgb <= "101111";
					when "010000010011001" => rgb <= "101111";
					when "010000010011010" => rgb <= "101111";
					when "010000010011011" => rgb <= "101111";
					when "010000010011100" => rgb <= "101111";
					when "010000010011101" => rgb <= "101111";
					when "010000010011110" => rgb <= "101111";
					when "010000010011111" => rgb <= "101111";
					when "010000100000000" => rgb <= "001000";
					when "010000100000001" => rgb <= "001000";
					when "010000100000010" => rgb <= "001000";
					when "010000100000011" => rgb <= "001000";
					when "010000100000100" => rgb <= "001000";
					when "010000100000101" => rgb <= "001000";
					when "010000100000110" => rgb <= "001000";
					when "010000100000111" => rgb <= "001000";
					when "010000100001000" => rgb <= "001000";
					when "010000100001001" => rgb <= "001000";
					when "010000100001010" => rgb <= "001000";
					when "010000100001011" => rgb <= "001000";
					when "010000100001100" => rgb <= "001000";
					when "010000100001101" => rgb <= "001000";
					when "010000100001110" => rgb <= "001000";
					when "010000100001111" => rgb <= "001000";
					when "010000100010000" => rgb <= "001000";
					when "010000100010001" => rgb <= "001000";
					when "010000100010010" => rgb <= "001000";
					when "010000100010011" => rgb <= "001000";
					when "010000100010100" => rgb <= "001000";
					when "010000100010101" => rgb <= "001000";
					when "010000100010110" => rgb <= "001000";
					when "010000100010111" => rgb <= "001000";
					when "010000100011000" => rgb <= "001000";
					when "010000100011001" => rgb <= "001000";
					when "010000100011010" => rgb <= "001000";
					when "010000100011011" => rgb <= "001000";
					when "010000100011100" => rgb <= "001000";
					when "010000100011101" => rgb <= "001000";
					when "010000100011110" => rgb <= "001000";
					when "010000100011111" => rgb <= "001000";
					when "010000100100000" => rgb <= "001000";
					when "010000100100001" => rgb <= "001000";
					when "010000100100010" => rgb <= "001000";
					when "010000100100011" => rgb <= "001000";
					when "010000100100100" => rgb <= "001000";
					when "010000100100101" => rgb <= "001000";
					when "010000100100110" => rgb <= "001000";
					when "010000100100111" => rgb <= "001000";
					when "010000100101000" => rgb <= "001000";
					when "010000100101001" => rgb <= "001000";
					when "010000100101010" => rgb <= "001000";
					when "010000100101011" => rgb <= "001000";
					when "010000100101100" => rgb <= "001000";
					when "010000100101101" => rgb <= "001000";
					when "010000100101110" => rgb <= "001000";
					when "010000100101111" => rgb <= "001000";
					when "010000100110000" => rgb <= "001000";
					when "010000100110001" => rgb <= "001000";
					when "010000100110010" => rgb <= "001000";
					when "010000100110011" => rgb <= "001000";
					when "010000100110100" => rgb <= "001000";
					when "010000100110101" => rgb <= "001000";
					when "010000100110110" => rgb <= "001000";
					when "010000100110111" => rgb <= "001000";
					when "010000100111000" => rgb <= "001000";
					when "010000100111001" => rgb <= "001000";
					when "010000100111010" => rgb <= "001000";
					when "010000100111011" => rgb <= "001000";
					when "010000100111100" => rgb <= "001000";
					when "010000100111101" => rgb <= "001000";
					when "010000100111110" => rgb <= "001000";
					when "010000100111111" => rgb <= "001000";
					when "010000101000000" => rgb <= "001000";
					when "010000101000001" => rgb <= "001000";
					when "010000101000010" => rgb <= "001000";
					when "010000101000011" => rgb <= "001000";
					when "010000101000100" => rgb <= "001000";
					when "010000101000101" => rgb <= "001000";
					when "010000101000110" => rgb <= "001000";
					when "010000101000111" => rgb <= "001000";
					when "010000101001000" => rgb <= "001000";
					when "010000101001001" => rgb <= "001000";
					when "010000101001010" => rgb <= "001000";
					when "010000101001011" => rgb <= "001000";
					when "010000101001100" => rgb <= "001000";
					when "010000101001101" => rgb <= "001000";
					when "010000101001110" => rgb <= "001000";
					when "010000101001111" => rgb <= "001000";
					when "010000101010000" => rgb <= "001000";
					when "010000101010001" => rgb <= "001000";
					when "010000101010010" => rgb <= "001000";
					when "010000101010011" => rgb <= "001000";
					when "010000101010100" => rgb <= "001000";
					when "010000101010101" => rgb <= "001000";
					when "010000101010110" => rgb <= "001000";
					when "010000101010111" => rgb <= "001000";
					when "010000101011000" => rgb <= "001000";
					when "010000101011001" => rgb <= "001000";
					when "010000101011010" => rgb <= "000000";
					when "010000101011011" => rgb <= "000000";
					when "010000101011100" => rgb <= "101111";
					when "010000101011101" => rgb <= "101111";
					when "010000101011110" => rgb <= "101111";
					when "010000101011111" => rgb <= "101111";
					when "010000101100000" => rgb <= "101111";
					when "010000101100001" => rgb <= "101111";
					when "010000101100010" => rgb <= "101111";
					when "010000101100011" => rgb <= "101111";
					when "010000101100100" => rgb <= "101111";
					when "010000101100101" => rgb <= "101111";
					when "010000101100110" => rgb <= "101111";
					when "010000101100111" => rgb <= "101111";
					when "010000101101000" => rgb <= "101111";
					when "010000101101001" => rgb <= "101111";
					when "010000101101010" => rgb <= "101111";
					when "010000101101011" => rgb <= "101111";
					when "010000101101100" => rgb <= "101111";
					when "010000101101101" => rgb <= "101111";
					when "010000101101110" => rgb <= "101111";
					when "010000101101111" => rgb <= "101111";
					when "010000101110000" => rgb <= "101111";
					when "010000101110001" => rgb <= "101111";
					when "010000101110010" => rgb <= "101111";
					when "010000101110011" => rgb <= "101111";
					when "010000101110100" => rgb <= "101111";
					when "010000101110101" => rgb <= "101111";
					when "010000101110110" => rgb <= "101111";
					when "010000101110111" => rgb <= "101111";
					when "010000101111000" => rgb <= "101111";
					when "010000101111001" => rgb <= "101111";
					when "010000101111010" => rgb <= "101111";
					when "010000101111011" => rgb <= "101111";
					when "010000101111100" => rgb <= "101111";
					when "010000101111101" => rgb <= "101111";
					when "010000101111110" => rgb <= "101111";
					when "010000101111111" => rgb <= "101111";
					when "010000110000000" => rgb <= "101111";
					when "010000110000001" => rgb <= "101111";
					when "010000110000010" => rgb <= "101111";
					when "010000110000011" => rgb <= "101111";
					when "010000110000100" => rgb <= "101111";
					when "010000110000101" => rgb <= "101111";
					when "010000110000110" => rgb <= "101111";
					when "010000110000111" => rgb <= "101111";
					when "010000110001000" => rgb <= "101111";
					when "010000110001001" => rgb <= "101111";
					when "010000110001010" => rgb <= "101111";
					when "010000110001011" => rgb <= "101111";
					when "010000110001100" => rgb <= "101111";
					when "010000110001101" => rgb <= "101111";
					when "010000110001110" => rgb <= "101111";
					when "010000110001111" => rgb <= "101111";
					when "010000110010000" => rgb <= "101111";
					when "010000110010001" => rgb <= "101111";
					when "010000110010010" => rgb <= "101111";
					when "010000110010011" => rgb <= "101111";
					when "010000110010100" => rgb <= "101111";
					when "010000110010101" => rgb <= "101111";
					when "010000110010110" => rgb <= "101111";
					when "010000110010111" => rgb <= "101111";
					when "010000110011000" => rgb <= "101111";
					when "010000110011001" => rgb <= "101111";
					when "010000110011010" => rgb <= "101111";
					when "010000110011011" => rgb <= "101111";
					when "010000110011100" => rgb <= "101111";
					when "010000110011101" => rgb <= "101111";
					when "010000110011110" => rgb <= "101111";
					when "010000110011111" => rgb <= "101111";
					when "010001000000000" => rgb <= "001000";
					when "010001000000001" => rgb <= "001000";
					when "010001000000010" => rgb <= "001000";
					when "010001000000011" => rgb <= "001000";
					when "010001000000100" => rgb <= "001000";
					when "010001000000101" => rgb <= "001000";
					when "010001000000110" => rgb <= "001000";
					when "010001000000111" => rgb <= "001000";
					when "010001000001000" => rgb <= "001000";
					when "010001000001001" => rgb <= "001000";
					when "010001000001010" => rgb <= "001000";
					when "010001000001011" => rgb <= "001000";
					when "010001000001100" => rgb <= "001000";
					when "010001000001101" => rgb <= "001000";
					when "010001000001110" => rgb <= "001000";
					when "010001000001111" => rgb <= "001000";
					when "010001000010000" => rgb <= "001000";
					when "010001000010001" => rgb <= "001000";
					when "010001000010010" => rgb <= "001000";
					when "010001000010011" => rgb <= "001000";
					when "010001000010100" => rgb <= "001000";
					when "010001000010101" => rgb <= "001000";
					when "010001000010110" => rgb <= "001000";
					when "010001000010111" => rgb <= "001000";
					when "010001000011000" => rgb <= "001000";
					when "010001000011001" => rgb <= "001000";
					when "010001000011010" => rgb <= "001000";
					when "010001000011011" => rgb <= "001000";
					when "010001000011100" => rgb <= "001000";
					when "010001000011101" => rgb <= "001000";
					when "010001000011110" => rgb <= "001000";
					when "010001000011111" => rgb <= "001000";
					when "010001000100000" => rgb <= "001000";
					when "010001000100001" => rgb <= "001000";
					when "010001000100010" => rgb <= "001000";
					when "010001000100011" => rgb <= "001000";
					when "010001000100100" => rgb <= "001000";
					when "010001000100101" => rgb <= "001000";
					when "010001000100110" => rgb <= "001000";
					when "010001000100111" => rgb <= "001000";
					when "010001000101000" => rgb <= "001000";
					when "010001000101001" => rgb <= "001000";
					when "010001000101010" => rgb <= "001000";
					when "010001000101011" => rgb <= "001000";
					when "010001000101100" => rgb <= "001000";
					when "010001000101101" => rgb <= "001000";
					when "010001000101110" => rgb <= "001000";
					when "010001000101111" => rgb <= "001000";
					when "010001000110000" => rgb <= "001000";
					when "010001000110001" => rgb <= "001000";
					when "010001000110010" => rgb <= "001000";
					when "010001000110011" => rgb <= "001000";
					when "010001000110100" => rgb <= "001000";
					when "010001000110101" => rgb <= "001000";
					when "010001000110110" => rgb <= "001000";
					when "010001000110111" => rgb <= "001000";
					when "010001000111000" => rgb <= "001000";
					when "010001000111001" => rgb <= "001000";
					when "010001000111010" => rgb <= "001000";
					when "010001000111011" => rgb <= "001000";
					when "010001000111100" => rgb <= "001000";
					when "010001000111101" => rgb <= "001000";
					when "010001000111110" => rgb <= "001000";
					when "010001000111111" => rgb <= "001000";
					when "010001001000000" => rgb <= "001000";
					when "010001001000001" => rgb <= "001000";
					when "010001001000010" => rgb <= "001000";
					when "010001001000011" => rgb <= "001000";
					when "010001001000100" => rgb <= "001000";
					when "010001001000101" => rgb <= "001000";
					when "010001001000110" => rgb <= "001000";
					when "010001001000111" => rgb <= "001000";
					when "010001001001000" => rgb <= "001000";
					when "010001001001001" => rgb <= "001000";
					when "010001001001010" => rgb <= "001000";
					when "010001001001011" => rgb <= "001000";
					when "010001001001100" => rgb <= "001000";
					when "010001001001101" => rgb <= "001000";
					when "010001001001110" => rgb <= "001000";
					when "010001001001111" => rgb <= "001000";
					when "010001001010000" => rgb <= "001000";
					when "010001001010001" => rgb <= "001000";
					when "010001001010010" => rgb <= "001000";
					when "010001001010011" => rgb <= "001000";
					when "010001001010100" => rgb <= "001000";
					when "010001001010101" => rgb <= "001000";
					when "010001001010110" => rgb <= "001000";
					when "010001001010111" => rgb <= "001000";
					when "010001001011000" => rgb <= "001000";
					when "010001001011001" => rgb <= "001000";
					when "010001001011010" => rgb <= "000000";
					when "010001001011011" => rgb <= "000000";
					when "010001001011100" => rgb <= "101111";
					when "010001001011101" => rgb <= "101111";
					when "010001001011110" => rgb <= "101111";
					when "010001001011111" => rgb <= "101111";
					when "010001001100000" => rgb <= "101111";
					when "010001001100001" => rgb <= "101111";
					when "010001001100010" => rgb <= "101111";
					when "010001001100011" => rgb <= "101111";
					when "010001001100100" => rgb <= "101111";
					when "010001001100101" => rgb <= "101111";
					when "010001001100110" => rgb <= "101111";
					when "010001001100111" => rgb <= "101111";
					when "010001001101000" => rgb <= "101111";
					when "010001001101001" => rgb <= "101111";
					when "010001001101010" => rgb <= "101111";
					when "010001001101011" => rgb <= "101111";
					when "010001001101100" => rgb <= "101111";
					when "010001001101101" => rgb <= "101111";
					when "010001001101110" => rgb <= "101111";
					when "010001001101111" => rgb <= "101111";
					when "010001001110000" => rgb <= "101111";
					when "010001001110001" => rgb <= "101111";
					when "010001001110010" => rgb <= "101111";
					when "010001001110011" => rgb <= "101111";
					when "010001001110100" => rgb <= "101111";
					when "010001001110101" => rgb <= "101111";
					when "010001001110110" => rgb <= "101111";
					when "010001001110111" => rgb <= "101111";
					when "010001001111000" => rgb <= "101111";
					when "010001001111001" => rgb <= "101111";
					when "010001001111010" => rgb <= "101111";
					when "010001001111011" => rgb <= "101111";
					when "010001001111100" => rgb <= "101111";
					when "010001001111101" => rgb <= "101111";
					when "010001001111110" => rgb <= "101111";
					when "010001001111111" => rgb <= "101111";
					when "010001010000000" => rgb <= "101111";
					when "010001010000001" => rgb <= "101111";
					when "010001010000010" => rgb <= "101111";
					when "010001010000011" => rgb <= "101111";
					when "010001010000100" => rgb <= "101111";
					when "010001010000101" => rgb <= "101111";
					when "010001010000110" => rgb <= "101111";
					when "010001010000111" => rgb <= "101111";
					when "010001010001000" => rgb <= "101111";
					when "010001010001001" => rgb <= "101111";
					when "010001010001010" => rgb <= "101111";
					when "010001010001011" => rgb <= "101111";
					when "010001010001100" => rgb <= "101111";
					when "010001010001101" => rgb <= "101111";
					when "010001010001110" => rgb <= "101111";
					when "010001010001111" => rgb <= "101111";
					when "010001010010000" => rgb <= "101111";
					when "010001010010001" => rgb <= "101111";
					when "010001010010010" => rgb <= "101111";
					when "010001010010011" => rgb <= "101111";
					when "010001010010100" => rgb <= "101111";
					when "010001010010101" => rgb <= "101111";
					when "010001010010110" => rgb <= "101111";
					when "010001010010111" => rgb <= "101111";
					when "010001010011000" => rgb <= "101111";
					when "010001010011001" => rgb <= "101111";
					when "010001010011010" => rgb <= "101111";
					when "010001010011011" => rgb <= "101111";
					when "010001010011100" => rgb <= "101111";
					when "010001010011101" => rgb <= "101111";
					when "010001010011110" => rgb <= "101111";
					when "010001010011111" => rgb <= "101111";
					when "010001100000000" => rgb <= "001000";
					when "010001100000001" => rgb <= "001000";
					when "010001100000010" => rgb <= "001000";
					when "010001100000011" => rgb <= "001000";
					when "010001100000100" => rgb <= "001000";
					when "010001100000101" => rgb <= "001000";
					when "010001100000110" => rgb <= "001000";
					when "010001100000111" => rgb <= "001000";
					when "010001100001000" => rgb <= "001000";
					when "010001100001001" => rgb <= "001000";
					when "010001100001010" => rgb <= "001000";
					when "010001100001011" => rgb <= "001000";
					when "010001100001100" => rgb <= "001000";
					when "010001100001101" => rgb <= "001000";
					when "010001100001110" => rgb <= "001000";
					when "010001100001111" => rgb <= "001000";
					when "010001100010000" => rgb <= "001000";
					when "010001100010001" => rgb <= "001000";
					when "010001100010010" => rgb <= "001000";
					when "010001100010011" => rgb <= "001000";
					when "010001100010100" => rgb <= "001000";
					when "010001100010101" => rgb <= "001000";
					when "010001100010110" => rgb <= "001000";
					when "010001100010111" => rgb <= "001000";
					when "010001100011000" => rgb <= "001000";
					when "010001100011001" => rgb <= "001000";
					when "010001100011010" => rgb <= "001000";
					when "010001100011011" => rgb <= "001000";
					when "010001100011100" => rgb <= "001000";
					when "010001100011101" => rgb <= "001000";
					when "010001100011110" => rgb <= "001000";
					when "010001100011111" => rgb <= "001000";
					when "010001100100000" => rgb <= "001000";
					when "010001100100001" => rgb <= "001000";
					when "010001100100010" => rgb <= "001000";
					when "010001100100011" => rgb <= "001000";
					when "010001100100100" => rgb <= "001000";
					when "010001100100101" => rgb <= "001000";
					when "010001100100110" => rgb <= "001000";
					when "010001100100111" => rgb <= "001000";
					when "010001100101000" => rgb <= "001000";
					when "010001100101001" => rgb <= "001000";
					when "010001100101010" => rgb <= "001000";
					when "010001100101011" => rgb <= "001000";
					when "010001100101100" => rgb <= "001000";
					when "010001100101101" => rgb <= "001000";
					when "010001100101110" => rgb <= "001000";
					when "010001100101111" => rgb <= "001000";
					when "010001100110000" => rgb <= "001000";
					when "010001100110001" => rgb <= "001000";
					when "010001100110010" => rgb <= "001000";
					when "010001100110011" => rgb <= "001000";
					when "010001100110100" => rgb <= "001000";
					when "010001100110101" => rgb <= "001000";
					when "010001100110110" => rgb <= "001000";
					when "010001100110111" => rgb <= "001000";
					when "010001100111000" => rgb <= "001000";
					when "010001100111001" => rgb <= "001000";
					when "010001100111010" => rgb <= "001000";
					when "010001100111011" => rgb <= "001000";
					when "010001100111100" => rgb <= "001000";
					when "010001100111101" => rgb <= "001000";
					when "010001100111110" => rgb <= "001000";
					when "010001100111111" => rgb <= "001000";
					when "010001101000000" => rgb <= "001000";
					when "010001101000001" => rgb <= "001000";
					when "010001101000010" => rgb <= "001000";
					when "010001101000011" => rgb <= "001000";
					when "010001101000100" => rgb <= "001000";
					when "010001101000101" => rgb <= "001000";
					when "010001101000110" => rgb <= "001000";
					when "010001101000111" => rgb <= "001000";
					when "010001101001000" => rgb <= "001000";
					when "010001101001001" => rgb <= "001000";
					when "010001101001010" => rgb <= "001000";
					when "010001101001011" => rgb <= "001000";
					when "010001101001100" => rgb <= "001000";
					when "010001101001101" => rgb <= "001000";
					when "010001101001110" => rgb <= "001000";
					when "010001101001111" => rgb <= "001000";
					when "010001101010000" => rgb <= "001000";
					when "010001101010001" => rgb <= "001000";
					when "010001101010010" => rgb <= "001000";
					when "010001101010011" => rgb <= "001000";
					when "010001101010100" => rgb <= "001000";
					when "010001101010101" => rgb <= "001000";
					when "010001101010110" => rgb <= "001000";
					when "010001101010111" => rgb <= "001000";
					when "010001101011000" => rgb <= "001000";
					when "010001101011001" => rgb <= "001000";
					when "010001101011010" => rgb <= "000000";
					when "010001101011011" => rgb <= "000000";
					when "010001101011100" => rgb <= "101111";
					when "010001101011101" => rgb <= "101111";
					when "010001101011110" => rgb <= "101111";
					when "010001101011111" => rgb <= "101111";
					when "010001101100000" => rgb <= "101111";
					when "010001101100001" => rgb <= "101111";
					when "010001101100010" => rgb <= "101111";
					when "010001101100011" => rgb <= "101111";
					when "010001101100100" => rgb <= "101111";
					when "010001101100101" => rgb <= "101111";
					when "010001101100110" => rgb <= "101111";
					when "010001101100111" => rgb <= "101111";
					when "010001101101000" => rgb <= "101111";
					when "010001101101001" => rgb <= "101111";
					when "010001101101010" => rgb <= "101111";
					when "010001101101011" => rgb <= "101111";
					when "010001101101100" => rgb <= "101111";
					when "010001101101101" => rgb <= "101111";
					when "010001101101110" => rgb <= "101111";
					when "010001101101111" => rgb <= "101111";
					when "010001101110000" => rgb <= "101111";
					when "010001101110001" => rgb <= "101111";
					when "010001101110010" => rgb <= "101111";
					when "010001101110011" => rgb <= "101111";
					when "010001101110100" => rgb <= "101111";
					when "010001101110101" => rgb <= "101111";
					when "010001101110110" => rgb <= "101111";
					when "010001101110111" => rgb <= "101111";
					when "010001101111000" => rgb <= "101111";
					when "010001101111001" => rgb <= "101111";
					when "010001101111010" => rgb <= "101111";
					when "010001101111011" => rgb <= "101111";
					when "010001101111100" => rgb <= "101111";
					when "010001101111101" => rgb <= "101111";
					when "010001101111110" => rgb <= "101111";
					when "010001101111111" => rgb <= "101111";
					when "010001110000000" => rgb <= "101111";
					when "010001110000001" => rgb <= "101111";
					when "010001110000010" => rgb <= "101111";
					when "010001110000011" => rgb <= "101111";
					when "010001110000100" => rgb <= "101111";
					when "010001110000101" => rgb <= "101111";
					when "010001110000110" => rgb <= "101111";
					when "010001110000111" => rgb <= "101111";
					when "010001110001000" => rgb <= "101111";
					when "010001110001001" => rgb <= "101111";
					when "010001110001010" => rgb <= "101111";
					when "010001110001011" => rgb <= "101111";
					when "010001110001100" => rgb <= "101111";
					when "010001110001101" => rgb <= "101111";
					when "010001110001110" => rgb <= "101111";
					when "010001110001111" => rgb <= "101111";
					when "010001110010000" => rgb <= "101111";
					when "010001110010001" => rgb <= "101111";
					when "010001110010010" => rgb <= "101111";
					when "010001110010011" => rgb <= "101111";
					when "010001110010100" => rgb <= "101111";
					when "010001110010101" => rgb <= "101111";
					when "010001110010110" => rgb <= "101111";
					when "010001110010111" => rgb <= "101111";
					when "010001110011000" => rgb <= "101111";
					when "010001110011001" => rgb <= "101111";
					when "010001110011010" => rgb <= "101111";
					when "010001110011011" => rgb <= "101111";
					when "010001110011100" => rgb <= "101111";
					when "010001110011101" => rgb <= "101111";
					when "010001110011110" => rgb <= "101111";
					when "010001110011111" => rgb <= "101111";
					when "010010000000000" => rgb <= "001000";
					when "010010000000001" => rgb <= "001000";
					when "010010000000010" => rgb <= "001000";
					when "010010000000011" => rgb <= "001000";
					when "010010000000100" => rgb <= "001000";
					when "010010000000101" => rgb <= "001000";
					when "010010000000110" => rgb <= "001000";
					when "010010000000111" => rgb <= "001000";
					when "010010000001000" => rgb <= "001000";
					when "010010000001001" => rgb <= "001000";
					when "010010000001010" => rgb <= "001000";
					when "010010000001011" => rgb <= "001000";
					when "010010000001100" => rgb <= "001000";
					when "010010000001101" => rgb <= "001000";
					when "010010000001110" => rgb <= "001000";
					when "010010000001111" => rgb <= "001000";
					when "010010000010000" => rgb <= "001000";
					when "010010000010001" => rgb <= "001000";
					when "010010000010010" => rgb <= "001000";
					when "010010000010011" => rgb <= "001000";
					when "010010000010100" => rgb <= "001000";
					when "010010000010101" => rgb <= "001000";
					when "010010000010110" => rgb <= "001000";
					when "010010000010111" => rgb <= "001000";
					when "010010000011000" => rgb <= "001000";
					when "010010000011001" => rgb <= "001000";
					when "010010000011010" => rgb <= "001000";
					when "010010000011011" => rgb <= "001000";
					when "010010000011100" => rgb <= "001000";
					when "010010000011101" => rgb <= "001000";
					when "010010000011110" => rgb <= "001000";
					when "010010000011111" => rgb <= "001000";
					when "010010000100000" => rgb <= "001000";
					when "010010000100001" => rgb <= "001000";
					when "010010000100010" => rgb <= "001000";
					when "010010000100011" => rgb <= "001000";
					when "010010000100100" => rgb <= "001000";
					when "010010000100101" => rgb <= "001000";
					when "010010000100110" => rgb <= "001000";
					when "010010000100111" => rgb <= "001000";
					when "010010000101000" => rgb <= "001000";
					when "010010000101001" => rgb <= "001000";
					when "010010000101010" => rgb <= "001000";
					when "010010000101011" => rgb <= "001000";
					when "010010000101100" => rgb <= "001000";
					when "010010000101101" => rgb <= "001000";
					when "010010000101110" => rgb <= "001000";
					when "010010000101111" => rgb <= "001000";
					when "010010000110000" => rgb <= "001000";
					when "010010000110001" => rgb <= "001000";
					when "010010000110010" => rgb <= "001000";
					when "010010000110011" => rgb <= "001000";
					when "010010000110100" => rgb <= "001000";
					when "010010000110101" => rgb <= "001000";
					when "010010000110110" => rgb <= "001000";
					when "010010000110111" => rgb <= "001000";
					when "010010000111000" => rgb <= "001000";
					when "010010000111001" => rgb <= "001000";
					when "010010000111010" => rgb <= "001000";
					when "010010000111011" => rgb <= "001000";
					when "010010000111100" => rgb <= "001000";
					when "010010000111101" => rgb <= "001000";
					when "010010000111110" => rgb <= "001000";
					when "010010000111111" => rgb <= "001000";
					when "010010001000000" => rgb <= "001000";
					when "010010001000001" => rgb <= "001000";
					when "010010001000010" => rgb <= "001000";
					when "010010001000011" => rgb <= "001000";
					when "010010001000100" => rgb <= "001000";
					when "010010001000101" => rgb <= "001000";
					when "010010001000110" => rgb <= "001000";
					when "010010001000111" => rgb <= "001000";
					when "010010001001000" => rgb <= "001000";
					when "010010001001001" => rgb <= "001000";
					when "010010001001010" => rgb <= "001000";
					when "010010001001011" => rgb <= "001000";
					when "010010001001100" => rgb <= "001000";
					when "010010001001101" => rgb <= "001000";
					when "010010001001110" => rgb <= "001000";
					when "010010001001111" => rgb <= "001000";
					when "010010001010000" => rgb <= "001000";
					when "010010001010001" => rgb <= "001000";
					when "010010001010010" => rgb <= "001000";
					when "010010001010011" => rgb <= "001000";
					when "010010001010100" => rgb <= "001000";
					when "010010001010101" => rgb <= "001000";
					when "010010001010110" => rgb <= "001000";
					when "010010001010111" => rgb <= "001000";
					when "010010001011000" => rgb <= "001000";
					when "010010001011001" => rgb <= "001000";
					when "010010001011010" => rgb <= "000000";
					when "010010001011011" => rgb <= "000000";
					when "010010001011100" => rgb <= "101111";
					when "010010001011101" => rgb <= "101111";
					when "010010001011110" => rgb <= "101111";
					when "010010001011111" => rgb <= "101111";
					when "010010001100000" => rgb <= "101111";
					when "010010001100001" => rgb <= "101111";
					when "010010001100010" => rgb <= "101111";
					when "010010001100011" => rgb <= "101111";
					when "010010001100100" => rgb <= "101111";
					when "010010001100101" => rgb <= "101111";
					when "010010001100110" => rgb <= "101111";
					when "010010001100111" => rgb <= "101111";
					when "010010001101000" => rgb <= "101111";
					when "010010001101001" => rgb <= "101111";
					when "010010001101010" => rgb <= "101111";
					when "010010001101011" => rgb <= "101111";
					when "010010001101100" => rgb <= "101111";
					when "010010001101101" => rgb <= "101111";
					when "010010001101110" => rgb <= "101111";
					when "010010001101111" => rgb <= "101111";
					when "010010001110000" => rgb <= "101111";
					when "010010001110001" => rgb <= "101111";
					when "010010001110010" => rgb <= "101111";
					when "010010001110011" => rgb <= "101111";
					when "010010001110100" => rgb <= "101111";
					when "010010001110101" => rgb <= "101111";
					when "010010001110110" => rgb <= "101111";
					when "010010001110111" => rgb <= "101111";
					when "010010001111000" => rgb <= "101111";
					when "010010001111001" => rgb <= "101111";
					when "010010001111010" => rgb <= "101111";
					when "010010001111011" => rgb <= "101111";
					when "010010001111100" => rgb <= "101111";
					when "010010001111101" => rgb <= "101111";
					when "010010001111110" => rgb <= "101111";
					when "010010001111111" => rgb <= "101111";
					when "010010010000000" => rgb <= "101111";
					when "010010010000001" => rgb <= "101111";
					when "010010010000010" => rgb <= "101111";
					when "010010010000011" => rgb <= "101111";
					when "010010010000100" => rgb <= "101111";
					when "010010010000101" => rgb <= "101111";
					when "010010010000110" => rgb <= "101111";
					when "010010010000111" => rgb <= "101111";
					when "010010010001000" => rgb <= "101111";
					when "010010010001001" => rgb <= "101111";
					when "010010010001010" => rgb <= "101111";
					when "010010010001011" => rgb <= "101111";
					when "010010010001100" => rgb <= "101111";
					when "010010010001101" => rgb <= "101111";
					when "010010010001110" => rgb <= "101111";
					when "010010010001111" => rgb <= "101111";
					when "010010010010000" => rgb <= "101111";
					when "010010010010001" => rgb <= "101111";
					when "010010010010010" => rgb <= "101111";
					when "010010010010011" => rgb <= "101111";
					when "010010010010100" => rgb <= "101111";
					when "010010010010101" => rgb <= "101111";
					when "010010010010110" => rgb <= "101111";
					when "010010010010111" => rgb <= "101111";
					when "010010010011000" => rgb <= "101111";
					when "010010010011001" => rgb <= "101111";
					when "010010010011010" => rgb <= "101111";
					when "010010010011011" => rgb <= "101111";
					when "010010010011100" => rgb <= "101111";
					when "010010010011101" => rgb <= "101111";
					when "010010010011110" => rgb <= "101111";
					when "010010010011111" => rgb <= "101111";
					when "010010100000000" => rgb <= "001000";
					when "010010100000001" => rgb <= "001000";
					when "010010100000010" => rgb <= "001000";
					when "010010100000011" => rgb <= "001000";
					when "010010100000100" => rgb <= "001000";
					when "010010100000101" => rgb <= "001000";
					when "010010100000110" => rgb <= "001000";
					when "010010100000111" => rgb <= "001000";
					when "010010100001000" => rgb <= "001000";
					when "010010100001001" => rgb <= "001000";
					when "010010100001010" => rgb <= "001000";
					when "010010100001011" => rgb <= "001000";
					when "010010100001100" => rgb <= "001000";
					when "010010100001101" => rgb <= "001000";
					when "010010100001110" => rgb <= "001000";
					when "010010100001111" => rgb <= "001000";
					when "010010100010000" => rgb <= "001000";
					when "010010100010001" => rgb <= "001000";
					when "010010100010010" => rgb <= "001000";
					when "010010100010011" => rgb <= "001000";
					when "010010100010100" => rgb <= "001000";
					when "010010100010101" => rgb <= "001000";
					when "010010100010110" => rgb <= "001000";
					when "010010100010111" => rgb <= "001000";
					when "010010100011000" => rgb <= "001000";
					when "010010100011001" => rgb <= "001000";
					when "010010100011010" => rgb <= "001000";
					when "010010100011011" => rgb <= "001000";
					when "010010100011100" => rgb <= "001000";
					when "010010100011101" => rgb <= "001000";
					when "010010100011110" => rgb <= "001000";
					when "010010100011111" => rgb <= "001000";
					when "010010100100000" => rgb <= "001000";
					when "010010100100001" => rgb <= "001000";
					when "010010100100010" => rgb <= "001000";
					when "010010100100011" => rgb <= "001000";
					when "010010100100100" => rgb <= "001000";
					when "010010100100101" => rgb <= "001000";
					when "010010100100110" => rgb <= "001000";
					when "010010100100111" => rgb <= "001000";
					when "010010100101000" => rgb <= "001000";
					when "010010100101001" => rgb <= "001000";
					when "010010100101010" => rgb <= "001000";
					when "010010100101011" => rgb <= "001000";
					when "010010100101100" => rgb <= "001000";
					when "010010100101101" => rgb <= "001000";
					when "010010100101110" => rgb <= "001000";
					when "010010100101111" => rgb <= "001000";
					when "010010100110000" => rgb <= "001000";
					when "010010100110001" => rgb <= "001000";
					when "010010100110010" => rgb <= "001000";
					when "010010100110011" => rgb <= "001000";
					when "010010100110100" => rgb <= "001000";
					when "010010100110101" => rgb <= "001000";
					when "010010100110110" => rgb <= "001000";
					when "010010100110111" => rgb <= "001000";
					when "010010100111000" => rgb <= "001000";
					when "010010100111001" => rgb <= "001000";
					when "010010100111010" => rgb <= "001000";
					when "010010100111011" => rgb <= "001000";
					when "010010100111100" => rgb <= "001000";
					when "010010100111101" => rgb <= "001000";
					when "010010100111110" => rgb <= "001000";
					when "010010100111111" => rgb <= "001000";
					when "010010101000000" => rgb <= "001000";
					when "010010101000001" => rgb <= "001000";
					when "010010101000010" => rgb <= "001000";
					when "010010101000011" => rgb <= "001000";
					when "010010101000100" => rgb <= "001000";
					when "010010101000101" => rgb <= "001000";
					when "010010101000110" => rgb <= "001000";
					when "010010101000111" => rgb <= "001000";
					when "010010101001000" => rgb <= "001000";
					when "010010101001001" => rgb <= "001000";
					when "010010101001010" => rgb <= "001000";
					when "010010101001011" => rgb <= "001000";
					when "010010101001100" => rgb <= "001000";
					when "010010101001101" => rgb <= "001000";
					when "010010101001110" => rgb <= "001000";
					when "010010101001111" => rgb <= "001000";
					when "010010101010000" => rgb <= "001000";
					when "010010101010001" => rgb <= "001000";
					when "010010101010010" => rgb <= "001000";
					when "010010101010011" => rgb <= "001000";
					when "010010101010100" => rgb <= "001000";
					when "010010101010101" => rgb <= "001000";
					when "010010101010110" => rgb <= "001000";
					when "010010101010111" => rgb <= "001000";
					when "010010101011000" => rgb <= "001000";
					when "010010101011001" => rgb <= "001000";
					when "010010101011010" => rgb <= "000000";
					when "010010101011011" => rgb <= "000000";
					when "010010101011100" => rgb <= "101111";
					when "010010101011101" => rgb <= "101111";
					when "010010101011110" => rgb <= "101111";
					when "010010101011111" => rgb <= "101111";
					when "010010101100000" => rgb <= "101111";
					when "010010101100001" => rgb <= "101111";
					when "010010101100010" => rgb <= "101111";
					when "010010101100011" => rgb <= "101111";
					when "010010101100100" => rgb <= "101111";
					when "010010101100101" => rgb <= "101111";
					when "010010101100110" => rgb <= "101111";
					when "010010101100111" => rgb <= "101111";
					when "010010101101000" => rgb <= "101111";
					when "010010101101001" => rgb <= "101111";
					when "010010101101010" => rgb <= "101111";
					when "010010101101011" => rgb <= "101111";
					when "010010101101100" => rgb <= "101111";
					when "010010101101101" => rgb <= "101111";
					when "010010101101110" => rgb <= "101111";
					when "010010101101111" => rgb <= "101111";
					when "010010101110000" => rgb <= "101111";
					when "010010101110001" => rgb <= "101111";
					when "010010101110010" => rgb <= "101111";
					when "010010101110011" => rgb <= "101111";
					when "010010101110100" => rgb <= "101111";
					when "010010101110101" => rgb <= "101111";
					when "010010101110110" => rgb <= "101111";
					when "010010101110111" => rgb <= "101111";
					when "010010101111000" => rgb <= "101111";
					when "010010101111001" => rgb <= "101111";
					when "010010101111010" => rgb <= "101111";
					when "010010101111011" => rgb <= "101111";
					when "010010101111100" => rgb <= "101111";
					when "010010101111101" => rgb <= "101111";
					when "010010101111110" => rgb <= "101111";
					when "010010101111111" => rgb <= "101111";
					when "010010110000000" => rgb <= "101111";
					when "010010110000001" => rgb <= "101111";
					when "010010110000010" => rgb <= "101111";
					when "010010110000011" => rgb <= "101111";
					when "010010110000100" => rgb <= "101111";
					when "010010110000101" => rgb <= "101111";
					when "010010110000110" => rgb <= "101111";
					when "010010110000111" => rgb <= "101111";
					when "010010110001000" => rgb <= "101111";
					when "010010110001001" => rgb <= "101111";
					when "010010110001010" => rgb <= "101111";
					when "010010110001011" => rgb <= "101111";
					when "010010110001100" => rgb <= "101111";
					when "010010110001101" => rgb <= "101111";
					when "010010110001110" => rgb <= "101111";
					when "010010110001111" => rgb <= "101111";
					when "010010110010000" => rgb <= "101111";
					when "010010110010001" => rgb <= "101111";
					when "010010110010010" => rgb <= "101111";
					when "010010110010011" => rgb <= "101111";
					when "010010110010100" => rgb <= "101111";
					when "010010110010101" => rgb <= "101111";
					when "010010110010110" => rgb <= "101111";
					when "010010110010111" => rgb <= "101111";
					when "010010110011000" => rgb <= "101111";
					when "010010110011001" => rgb <= "101111";
					when "010010110011010" => rgb <= "101111";
					when "010010110011011" => rgb <= "101111";
					when "010010110011100" => rgb <= "101111";
					when "010010110011101" => rgb <= "101111";
					when "010010110011110" => rgb <= "101111";
					when "010010110011111" => rgb <= "101111";
					when "010011000000000" => rgb <= "001000";
					when "010011000000001" => rgb <= "001000";
					when "010011000000010" => rgb <= "001000";
					when "010011000000011" => rgb <= "001000";
					when "010011000000100" => rgb <= "001000";
					when "010011000000101" => rgb <= "001000";
					when "010011000000110" => rgb <= "001000";
					when "010011000000111" => rgb <= "001000";
					when "010011000001000" => rgb <= "001000";
					when "010011000001001" => rgb <= "001000";
					when "010011000001010" => rgb <= "001000";
					when "010011000001011" => rgb <= "001000";
					when "010011000001100" => rgb <= "001000";
					when "010011000001101" => rgb <= "001000";
					when "010011000001110" => rgb <= "001000";
					when "010011000001111" => rgb <= "001000";
					when "010011000010000" => rgb <= "001000";
					when "010011000010001" => rgb <= "001000";
					when "010011000010010" => rgb <= "001000";
					when "010011000010011" => rgb <= "001000";
					when "010011000010100" => rgb <= "001000";
					when "010011000010101" => rgb <= "001000";
					when "010011000010110" => rgb <= "001000";
					when "010011000010111" => rgb <= "001000";
					when "010011000011000" => rgb <= "001000";
					when "010011000011001" => rgb <= "001000";
					when "010011000011010" => rgb <= "001000";
					when "010011000011011" => rgb <= "001000";
					when "010011000011100" => rgb <= "001000";
					when "010011000011101" => rgb <= "001000";
					when "010011000011110" => rgb <= "001000";
					when "010011000011111" => rgb <= "001000";
					when "010011000100000" => rgb <= "001000";
					when "010011000100001" => rgb <= "001000";
					when "010011000100010" => rgb <= "001000";
					when "010011000100011" => rgb <= "001000";
					when "010011000100100" => rgb <= "001000";
					when "010011000100101" => rgb <= "001000";
					when "010011000100110" => rgb <= "001000";
					when "010011000100111" => rgb <= "001000";
					when "010011000101000" => rgb <= "001000";
					when "010011000101001" => rgb <= "001000";
					when "010011000101010" => rgb <= "001000";
					when "010011000101011" => rgb <= "001000";
					when "010011000101100" => rgb <= "001000";
					when "010011000101101" => rgb <= "001000";
					when "010011000101110" => rgb <= "001000";
					when "010011000101111" => rgb <= "001000";
					when "010011000110000" => rgb <= "001000";
					when "010011000110001" => rgb <= "001000";
					when "010011000110010" => rgb <= "001000";
					when "010011000110011" => rgb <= "001000";
					when "010011000110100" => rgb <= "001000";
					when "010011000110101" => rgb <= "001000";
					when "010011000110110" => rgb <= "001000";
					when "010011000110111" => rgb <= "001000";
					when "010011000111000" => rgb <= "001000";
					when "010011000111001" => rgb <= "001000";
					when "010011000111010" => rgb <= "001000";
					when "010011000111011" => rgb <= "001000";
					when "010011000111100" => rgb <= "001000";
					when "010011000111101" => rgb <= "001000";
					when "010011000111110" => rgb <= "001000";
					when "010011000111111" => rgb <= "001000";
					when "010011001000000" => rgb <= "001000";
					when "010011001000001" => rgb <= "001000";
					when "010011001000010" => rgb <= "001000";
					when "010011001000011" => rgb <= "001000";
					when "010011001000100" => rgb <= "001000";
					when "010011001000101" => rgb <= "001000";
					when "010011001000110" => rgb <= "001000";
					when "010011001000111" => rgb <= "001000";
					when "010011001001000" => rgb <= "001000";
					when "010011001001001" => rgb <= "001000";
					when "010011001001010" => rgb <= "001000";
					when "010011001001011" => rgb <= "001000";
					when "010011001001100" => rgb <= "001000";
					when "010011001001101" => rgb <= "001000";
					when "010011001001110" => rgb <= "001000";
					when "010011001001111" => rgb <= "001000";
					when "010011001010000" => rgb <= "001000";
					when "010011001010001" => rgb <= "001000";
					when "010011001010010" => rgb <= "001000";
					when "010011001010011" => rgb <= "001000";
					when "010011001010100" => rgb <= "001000";
					when "010011001010101" => rgb <= "001000";
					when "010011001010110" => rgb <= "001000";
					when "010011001010111" => rgb <= "001000";
					when "010011001011000" => rgb <= "001000";
					when "010011001011001" => rgb <= "001000";
					when "010011001011010" => rgb <= "000000";
					when "010011001011011" => rgb <= "000000";
					when "010011001011100" => rgb <= "101111";
					when "010011001011101" => rgb <= "101111";
					when "010011001011110" => rgb <= "101111";
					when "010011001011111" => rgb <= "101111";
					when "010011001100000" => rgb <= "101111";
					when "010011001100001" => rgb <= "101111";
					when "010011001100010" => rgb <= "101111";
					when "010011001100011" => rgb <= "101111";
					when "010011001100100" => rgb <= "101111";
					when "010011001100101" => rgb <= "101111";
					when "010011001100110" => rgb <= "101111";
					when "010011001100111" => rgb <= "101111";
					when "010011001101000" => rgb <= "101111";
					when "010011001101001" => rgb <= "101111";
					when "010011001101010" => rgb <= "101111";
					when "010011001101011" => rgb <= "101111";
					when "010011001101100" => rgb <= "101111";
					when "010011001101101" => rgb <= "101111";
					when "010011001101110" => rgb <= "101111";
					when "010011001101111" => rgb <= "101111";
					when "010011001110000" => rgb <= "101111";
					when "010011001110001" => rgb <= "101111";
					when "010011001110010" => rgb <= "101111";
					when "010011001110011" => rgb <= "101111";
					when "010011001110100" => rgb <= "101111";
					when "010011001110101" => rgb <= "101111";
					when "010011001110110" => rgb <= "101111";
					when "010011001110111" => rgb <= "101111";
					when "010011001111000" => rgb <= "101111";
					when "010011001111001" => rgb <= "101111";
					when "010011001111010" => rgb <= "101111";
					when "010011001111011" => rgb <= "101111";
					when "010011001111100" => rgb <= "101111";
					when "010011001111101" => rgb <= "101111";
					when "010011001111110" => rgb <= "101111";
					when "010011001111111" => rgb <= "101111";
					when "010011010000000" => rgb <= "101111";
					when "010011010000001" => rgb <= "101111";
					when "010011010000010" => rgb <= "101111";
					when "010011010000011" => rgb <= "101111";
					when "010011010000100" => rgb <= "101111";
					when "010011010000101" => rgb <= "101111";
					when "010011010000110" => rgb <= "101111";
					when "010011010000111" => rgb <= "101111";
					when "010011010001000" => rgb <= "101111";
					when "010011010001001" => rgb <= "101111";
					when "010011010001010" => rgb <= "101111";
					when "010011010001011" => rgb <= "101111";
					when "010011010001100" => rgb <= "101111";
					when "010011010001101" => rgb <= "101111";
					when "010011010001110" => rgb <= "101111";
					when "010011010001111" => rgb <= "101111";
					when "010011010010000" => rgb <= "101111";
					when "010011010010001" => rgb <= "101111";
					when "010011010010010" => rgb <= "101111";
					when "010011010010011" => rgb <= "101111";
					when "010011010010100" => rgb <= "101111";
					when "010011010010101" => rgb <= "101111";
					when "010011010010110" => rgb <= "101111";
					when "010011010010111" => rgb <= "101111";
					when "010011010011000" => rgb <= "101111";
					when "010011010011001" => rgb <= "101111";
					when "010011010011010" => rgb <= "101111";
					when "010011010011011" => rgb <= "101111";
					when "010011010011100" => rgb <= "101111";
					when "010011010011101" => rgb <= "101111";
					when "010011010011110" => rgb <= "101111";
					when "010011010011111" => rgb <= "101111";
					when "010011100000000" => rgb <= "001000";
					when "010011100000001" => rgb <= "001000";
					when "010011100000010" => rgb <= "001000";
					when "010011100000011" => rgb <= "001000";
					when "010011100000100" => rgb <= "001000";
					when "010011100000101" => rgb <= "001000";
					when "010011100000110" => rgb <= "001000";
					when "010011100000111" => rgb <= "001000";
					when "010011100001000" => rgb <= "001000";
					when "010011100001001" => rgb <= "001000";
					when "010011100001010" => rgb <= "001000";
					when "010011100001011" => rgb <= "001000";
					when "010011100001100" => rgb <= "001000";
					when "010011100001101" => rgb <= "001000";
					when "010011100001110" => rgb <= "001000";
					when "010011100001111" => rgb <= "001000";
					when "010011100010000" => rgb <= "001000";
					when "010011100010001" => rgb <= "001000";
					when "010011100010010" => rgb <= "001000";
					when "010011100010011" => rgb <= "001000";
					when "010011100010100" => rgb <= "001000";
					when "010011100010101" => rgb <= "001000";
					when "010011100010110" => rgb <= "001000";
					when "010011100010111" => rgb <= "001000";
					when "010011100011000" => rgb <= "001000";
					when "010011100011001" => rgb <= "001000";
					when "010011100011010" => rgb <= "001000";
					when "010011100011011" => rgb <= "001000";
					when "010011100011100" => rgb <= "001000";
					when "010011100011101" => rgb <= "001000";
					when "010011100011110" => rgb <= "001000";
					when "010011100011111" => rgb <= "001000";
					when "010011100100000" => rgb <= "001000";
					when "010011100100001" => rgb <= "001000";
					when "010011100100010" => rgb <= "001000";
					when "010011100100011" => rgb <= "001000";
					when "010011100100100" => rgb <= "001000";
					when "010011100100101" => rgb <= "001000";
					when "010011100100110" => rgb <= "001000";
					when "010011100100111" => rgb <= "001000";
					when "010011100101000" => rgb <= "001000";
					when "010011100101001" => rgb <= "001000";
					when "010011100101010" => rgb <= "001000";
					when "010011100101011" => rgb <= "001000";
					when "010011100101100" => rgb <= "001000";
					when "010011100101101" => rgb <= "001000";
					when "010011100101110" => rgb <= "001000";
					when "010011100101111" => rgb <= "001000";
					when "010011100110000" => rgb <= "001000";
					when "010011100110001" => rgb <= "001000";
					when "010011100110010" => rgb <= "001000";
					when "010011100110011" => rgb <= "001000";
					when "010011100110100" => rgb <= "001000";
					when "010011100110101" => rgb <= "001000";
					when "010011100110110" => rgb <= "001000";
					when "010011100110111" => rgb <= "001000";
					when "010011100111000" => rgb <= "001000";
					when "010011100111001" => rgb <= "001000";
					when "010011100111010" => rgb <= "001000";
					when "010011100111011" => rgb <= "001000";
					when "010011100111100" => rgb <= "001000";
					when "010011100111101" => rgb <= "001000";
					when "010011100111110" => rgb <= "001000";
					when "010011100111111" => rgb <= "001000";
					when "010011101000000" => rgb <= "001000";
					when "010011101000001" => rgb <= "001000";
					when "010011101000010" => rgb <= "001000";
					when "010011101000011" => rgb <= "001000";
					when "010011101000100" => rgb <= "001000";
					when "010011101000101" => rgb <= "001000";
					when "010011101000110" => rgb <= "001000";
					when "010011101000111" => rgb <= "001000";
					when "010011101001000" => rgb <= "001000";
					when "010011101001001" => rgb <= "001000";
					when "010011101001010" => rgb <= "001000";
					when "010011101001011" => rgb <= "001000";
					when "010011101001100" => rgb <= "001000";
					when "010011101001101" => rgb <= "001000";
					when "010011101001110" => rgb <= "001000";
					when "010011101001111" => rgb <= "001000";
					when "010011101010000" => rgb <= "001000";
					when "010011101010001" => rgb <= "001000";
					when "010011101010010" => rgb <= "001000";
					when "010011101010011" => rgb <= "001000";
					when "010011101010100" => rgb <= "001000";
					when "010011101010101" => rgb <= "001000";
					when "010011101010110" => rgb <= "001000";
					when "010011101010111" => rgb <= "001000";
					when "010011101011000" => rgb <= "001000";
					when "010011101011001" => rgb <= "001000";
					when "010011101011010" => rgb <= "000000";
					when "010011101011011" => rgb <= "000000";
					when "010011101011100" => rgb <= "101111";
					when "010011101011101" => rgb <= "101111";
					when "010011101011110" => rgb <= "101111";
					when "010011101011111" => rgb <= "101111";
					when "010011101100000" => rgb <= "101111";
					when "010011101100001" => rgb <= "101111";
					when "010011101100010" => rgb <= "101111";
					when "010011101100011" => rgb <= "101111";
					when "010011101100100" => rgb <= "101111";
					when "010011101100101" => rgb <= "101111";
					when "010011101100110" => rgb <= "101111";
					when "010011101100111" => rgb <= "101111";
					when "010011101101000" => rgb <= "101111";
					when "010011101101001" => rgb <= "101111";
					when "010011101101010" => rgb <= "101111";
					when "010011101101011" => rgb <= "101111";
					when "010011101101100" => rgb <= "101111";
					when "010011101101101" => rgb <= "101111";
					when "010011101101110" => rgb <= "101111";
					when "010011101101111" => rgb <= "101111";
					when "010011101110000" => rgb <= "101111";
					when "010011101110001" => rgb <= "101111";
					when "010011101110010" => rgb <= "101111";
					when "010011101110011" => rgb <= "101111";
					when "010011101110100" => rgb <= "101111";
					when "010011101110101" => rgb <= "101111";
					when "010011101110110" => rgb <= "101111";
					when "010011101110111" => rgb <= "101111";
					when "010011101111000" => rgb <= "101111";
					when "010011101111001" => rgb <= "101111";
					when "010011101111010" => rgb <= "101111";
					when "010011101111011" => rgb <= "101111";
					when "010011101111100" => rgb <= "101111";
					when "010011101111101" => rgb <= "101111";
					when "010011101111110" => rgb <= "101111";
					when "010011101111111" => rgb <= "101111";
					when "010011110000000" => rgb <= "101111";
					when "010011110000001" => rgb <= "101111";
					when "010011110000010" => rgb <= "101111";
					when "010011110000011" => rgb <= "101111";
					when "010011110000100" => rgb <= "101111";
					when "010011110000101" => rgb <= "101111";
					when "010011110000110" => rgb <= "101111";
					when "010011110000111" => rgb <= "101111";
					when "010011110001000" => rgb <= "101111";
					when "010011110001001" => rgb <= "101111";
					when "010011110001010" => rgb <= "101111";
					when "010011110001011" => rgb <= "101111";
					when "010011110001100" => rgb <= "101111";
					when "010011110001101" => rgb <= "101111";
					when "010011110001110" => rgb <= "101111";
					when "010011110001111" => rgb <= "101111";
					when "010011110010000" => rgb <= "101111";
					when "010011110010001" => rgb <= "101111";
					when "010011110010010" => rgb <= "101111";
					when "010011110010011" => rgb <= "101111";
					when "010011110010100" => rgb <= "101111";
					when "010011110010101" => rgb <= "101111";
					when "010011110010110" => rgb <= "101111";
					when "010011110010111" => rgb <= "101111";
					when "010011110011000" => rgb <= "101111";
					when "010011110011001" => rgb <= "101111";
					when "010011110011010" => rgb <= "101111";
					when "010011110011011" => rgb <= "101111";
					when "010011110011100" => rgb <= "101111";
					when "010011110011101" => rgb <= "101111";
					when "010011110011110" => rgb <= "101111";
					when "010011110011111" => rgb <= "101111";
					when "010100000000000" => rgb <= "001000";
					when "010100000000001" => rgb <= "001000";
					when "010100000000010" => rgb <= "001000";
					when "010100000000011" => rgb <= "001000";
					when "010100000000100" => rgb <= "001000";
					when "010100000000101" => rgb <= "001000";
					when "010100000000110" => rgb <= "001000";
					when "010100000000111" => rgb <= "001000";
					when "010100000001000" => rgb <= "001000";
					when "010100000001001" => rgb <= "001000";
					when "010100000001010" => rgb <= "001000";
					when "010100000001011" => rgb <= "001000";
					when "010100000001100" => rgb <= "001000";
					when "010100000001101" => rgb <= "001000";
					when "010100000001110" => rgb <= "001000";
					when "010100000001111" => rgb <= "001000";
					when "010100000010000" => rgb <= "001000";
					when "010100000010001" => rgb <= "001000";
					when "010100000010010" => rgb <= "001000";
					when "010100000010011" => rgb <= "001000";
					when "010100000010100" => rgb <= "001000";
					when "010100000010101" => rgb <= "001000";
					when "010100000010110" => rgb <= "001000";
					when "010100000010111" => rgb <= "001000";
					when "010100000011000" => rgb <= "001000";
					when "010100000011001" => rgb <= "001000";
					when "010100000011010" => rgb <= "001000";
					when "010100000011011" => rgb <= "001000";
					when "010100000011100" => rgb <= "001000";
					when "010100000011101" => rgb <= "001000";
					when "010100000011110" => rgb <= "001000";
					when "010100000011111" => rgb <= "001000";
					when "010100000100000" => rgb <= "001000";
					when "010100000100001" => rgb <= "001000";
					when "010100000100010" => rgb <= "001000";
					when "010100000100011" => rgb <= "001000";
					when "010100000100100" => rgb <= "001000";
					when "010100000100101" => rgb <= "001000";
					when "010100000100110" => rgb <= "001000";
					when "010100000100111" => rgb <= "001000";
					when "010100000101000" => rgb <= "001000";
					when "010100000101001" => rgb <= "001000";
					when "010100000101010" => rgb <= "001000";
					when "010100000101011" => rgb <= "001000";
					when "010100000101100" => rgb <= "001000";
					when "010100000101101" => rgb <= "001000";
					when "010100000101110" => rgb <= "001000";
					when "010100000101111" => rgb <= "001000";
					when "010100000110000" => rgb <= "001000";
					when "010100000110001" => rgb <= "001000";
					when "010100000110010" => rgb <= "001000";
					when "010100000110011" => rgb <= "001000";
					when "010100000110100" => rgb <= "001000";
					when "010100000110101" => rgb <= "001000";
					when "010100000110110" => rgb <= "001000";
					when "010100000110111" => rgb <= "001000";
					when "010100000111000" => rgb <= "001000";
					when "010100000111001" => rgb <= "001000";
					when "010100000111010" => rgb <= "001000";
					when "010100000111011" => rgb <= "001000";
					when "010100000111100" => rgb <= "001000";
					when "010100000111101" => rgb <= "001000";
					when "010100000111110" => rgb <= "001000";
					when "010100000111111" => rgb <= "001000";
					when "010100001000000" => rgb <= "001000";
					when "010100001000001" => rgb <= "001000";
					when "010100001000010" => rgb <= "001000";
					when "010100001000011" => rgb <= "001000";
					when "010100001000100" => rgb <= "001000";
					when "010100001000101" => rgb <= "001000";
					when "010100001000110" => rgb <= "001000";
					when "010100001000111" => rgb <= "001000";
					when "010100001001000" => rgb <= "001000";
					when "010100001001001" => rgb <= "001000";
					when "010100001001010" => rgb <= "001000";
					when "010100001001011" => rgb <= "001000";
					when "010100001001100" => rgb <= "001000";
					when "010100001001101" => rgb <= "001000";
					when "010100001001110" => rgb <= "001000";
					when "010100001001111" => rgb <= "001000";
					when "010100001010000" => rgb <= "001000";
					when "010100001010001" => rgb <= "001000";
					when "010100001010010" => rgb <= "001000";
					when "010100001010011" => rgb <= "001000";
					when "010100001010100" => rgb <= "001000";
					when "010100001010101" => rgb <= "001000";
					when "010100001010110" => rgb <= "001000";
					when "010100001010111" => rgb <= "001000";
					when "010100001011000" => rgb <= "000000";
					when "010100001011001" => rgb <= "000000";
					when "010100001011010" => rgb <= "000000";
					when "010100001011011" => rgb <= "000000";
					when "010100001011100" => rgb <= "101111";
					when "010100001011101" => rgb <= "101111";
					when "010100001011110" => rgb <= "101111";
					when "010100001011111" => rgb <= "101111";
					when "010100001100000" => rgb <= "101111";
					when "010100001100001" => rgb <= "101111";
					when "010100001100010" => rgb <= "101111";
					when "010100001100011" => rgb <= "101111";
					when "010100001100100" => rgb <= "101111";
					when "010100001100101" => rgb <= "101111";
					when "010100001100110" => rgb <= "101111";
					when "010100001100111" => rgb <= "101111";
					when "010100001101000" => rgb <= "101111";
					when "010100001101001" => rgb <= "101111";
					when "010100001101010" => rgb <= "101111";
					when "010100001101011" => rgb <= "101111";
					when "010100001101100" => rgb <= "101111";
					when "010100001101101" => rgb <= "101111";
					when "010100001101110" => rgb <= "101111";
					when "010100001101111" => rgb <= "101111";
					when "010100001110000" => rgb <= "101111";
					when "010100001110001" => rgb <= "101111";
					when "010100001110010" => rgb <= "101111";
					when "010100001110011" => rgb <= "101111";
					when "010100001110100" => rgb <= "101111";
					when "010100001110101" => rgb <= "101111";
					when "010100001110110" => rgb <= "101111";
					when "010100001110111" => rgb <= "101111";
					when "010100001111000" => rgb <= "101111";
					when "010100001111001" => rgb <= "101111";
					when "010100001111010" => rgb <= "101111";
					when "010100001111011" => rgb <= "101111";
					when "010100001111100" => rgb <= "101111";
					when "010100001111101" => rgb <= "101111";
					when "010100001111110" => rgb <= "101111";
					when "010100001111111" => rgb <= "101111";
					when "010100010000000" => rgb <= "101111";
					when "010100010000001" => rgb <= "101111";
					when "010100010000010" => rgb <= "101111";
					when "010100010000011" => rgb <= "101111";
					when "010100010000100" => rgb <= "101111";
					when "010100010000101" => rgb <= "101111";
					when "010100010000110" => rgb <= "101111";
					when "010100010000111" => rgb <= "101111";
					when "010100010001000" => rgb <= "101111";
					when "010100010001001" => rgb <= "101111";
					when "010100010001010" => rgb <= "101111";
					when "010100010001011" => rgb <= "101111";
					when "010100010001100" => rgb <= "101111";
					when "010100010001101" => rgb <= "101111";
					when "010100010001110" => rgb <= "101111";
					when "010100010001111" => rgb <= "101111";
					when "010100010010000" => rgb <= "101111";
					when "010100010010001" => rgb <= "101111";
					when "010100010010010" => rgb <= "101111";
					when "010100010010011" => rgb <= "101111";
					when "010100010010100" => rgb <= "101111";
					when "010100010010101" => rgb <= "101111";
					when "010100010010110" => rgb <= "101111";
					when "010100010010111" => rgb <= "101111";
					when "010100010011000" => rgb <= "101111";
					when "010100010011001" => rgb <= "101111";
					when "010100010011010" => rgb <= "101111";
					when "010100010011011" => rgb <= "101111";
					when "010100010011100" => rgb <= "101111";
					when "010100010011101" => rgb <= "101111";
					when "010100010011110" => rgb <= "101111";
					when "010100010011111" => rgb <= "101111";
					when "010100100000000" => rgb <= "001000";
					when "010100100000001" => rgb <= "001000";
					when "010100100000010" => rgb <= "001000";
					when "010100100000011" => rgb <= "001000";
					when "010100100000100" => rgb <= "001000";
					when "010100100000101" => rgb <= "001000";
					when "010100100000110" => rgb <= "001000";
					when "010100100000111" => rgb <= "001000";
					when "010100100001000" => rgb <= "001000";
					when "010100100001001" => rgb <= "001000";
					when "010100100001010" => rgb <= "001000";
					when "010100100001011" => rgb <= "001000";
					when "010100100001100" => rgb <= "001000";
					when "010100100001101" => rgb <= "001000";
					when "010100100001110" => rgb <= "001000";
					when "010100100001111" => rgb <= "001000";
					when "010100100010000" => rgb <= "001000";
					when "010100100010001" => rgb <= "001000";
					when "010100100010010" => rgb <= "001000";
					when "010100100010011" => rgb <= "001000";
					when "010100100010100" => rgb <= "001000";
					when "010100100010101" => rgb <= "001000";
					when "010100100010110" => rgb <= "001000";
					when "010100100010111" => rgb <= "001000";
					when "010100100011000" => rgb <= "001000";
					when "010100100011001" => rgb <= "001000";
					when "010100100011010" => rgb <= "001000";
					when "010100100011011" => rgb <= "001000";
					when "010100100011100" => rgb <= "001000";
					when "010100100011101" => rgb <= "001000";
					when "010100100011110" => rgb <= "001000";
					when "010100100011111" => rgb <= "001000";
					when "010100100100000" => rgb <= "001000";
					when "010100100100001" => rgb <= "001000";
					when "010100100100010" => rgb <= "001000";
					when "010100100100011" => rgb <= "001000";
					when "010100100100100" => rgb <= "001000";
					when "010100100100101" => rgb <= "001000";
					when "010100100100110" => rgb <= "001000";
					when "010100100100111" => rgb <= "001000";
					when "010100100101000" => rgb <= "001000";
					when "010100100101001" => rgb <= "001000";
					when "010100100101010" => rgb <= "001000";
					when "010100100101011" => rgb <= "001000";
					when "010100100101100" => rgb <= "001000";
					when "010100100101101" => rgb <= "001000";
					when "010100100101110" => rgb <= "001000";
					when "010100100101111" => rgb <= "001000";
					when "010100100110000" => rgb <= "001000";
					when "010100100110001" => rgb <= "001000";
					when "010100100110010" => rgb <= "001000";
					when "010100100110011" => rgb <= "001000";
					when "010100100110100" => rgb <= "001000";
					when "010100100110101" => rgb <= "001000";
					when "010100100110110" => rgb <= "001000";
					when "010100100110111" => rgb <= "001000";
					when "010100100111000" => rgb <= "001000";
					when "010100100111001" => rgb <= "001000";
					when "010100100111010" => rgb <= "001000";
					when "010100100111011" => rgb <= "001000";
					when "010100100111100" => rgb <= "001000";
					when "010100100111101" => rgb <= "001000";
					when "010100100111110" => rgb <= "001000";
					when "010100100111111" => rgb <= "001000";
					when "010100101000000" => rgb <= "001000";
					when "010100101000001" => rgb <= "001000";
					when "010100101000010" => rgb <= "001000";
					when "010100101000011" => rgb <= "001000";
					when "010100101000100" => rgb <= "001000";
					when "010100101000101" => rgb <= "001000";
					when "010100101000110" => rgb <= "001000";
					when "010100101000111" => rgb <= "001000";
					when "010100101001000" => rgb <= "001000";
					when "010100101001001" => rgb <= "001000";
					when "010100101001010" => rgb <= "001000";
					when "010100101001011" => rgb <= "001000";
					when "010100101001100" => rgb <= "001000";
					when "010100101001101" => rgb <= "001000";
					when "010100101001110" => rgb <= "001000";
					when "010100101001111" => rgb <= "001000";
					when "010100101010000" => rgb <= "001000";
					when "010100101010001" => rgb <= "001000";
					when "010100101010010" => rgb <= "001000";
					when "010100101010011" => rgb <= "001000";
					when "010100101010100" => rgb <= "001000";
					when "010100101010101" => rgb <= "001000";
					when "010100101010110" => rgb <= "001000";
					when "010100101010111" => rgb <= "001000";
					when "010100101011000" => rgb <= "000000";
					when "010100101011001" => rgb <= "000000";
					when "010100101011010" => rgb <= "000000";
					when "010100101011011" => rgb <= "000000";
					when "010100101011100" => rgb <= "101111";
					when "010100101011101" => rgb <= "101111";
					when "010100101011110" => rgb <= "101111";
					when "010100101011111" => rgb <= "101111";
					when "010100101100000" => rgb <= "101111";
					when "010100101100001" => rgb <= "101111";
					when "010100101100010" => rgb <= "101111";
					when "010100101100011" => rgb <= "101111";
					when "010100101100100" => rgb <= "101111";
					when "010100101100101" => rgb <= "101111";
					when "010100101100110" => rgb <= "101111";
					when "010100101100111" => rgb <= "101111";
					when "010100101101000" => rgb <= "101111";
					when "010100101101001" => rgb <= "101111";
					when "010100101101010" => rgb <= "101111";
					when "010100101101011" => rgb <= "101111";
					when "010100101101100" => rgb <= "101111";
					when "010100101101101" => rgb <= "101111";
					when "010100101101110" => rgb <= "101111";
					when "010100101101111" => rgb <= "101111";
					when "010100101110000" => rgb <= "101111";
					when "010100101110001" => rgb <= "101111";
					when "010100101110010" => rgb <= "101111";
					when "010100101110011" => rgb <= "101111";
					when "010100101110100" => rgb <= "101111";
					when "010100101110101" => rgb <= "101111";
					when "010100101110110" => rgb <= "101111";
					when "010100101110111" => rgb <= "101111";
					when "010100101111000" => rgb <= "101111";
					when "010100101111001" => rgb <= "101111";
					when "010100101111010" => rgb <= "101111";
					when "010100101111011" => rgb <= "101111";
					when "010100101111100" => rgb <= "101111";
					when "010100101111101" => rgb <= "101111";
					when "010100101111110" => rgb <= "101111";
					when "010100101111111" => rgb <= "101111";
					when "010100110000000" => rgb <= "101111";
					when "010100110000001" => rgb <= "101111";
					when "010100110000010" => rgb <= "101111";
					when "010100110000011" => rgb <= "101111";
					when "010100110000100" => rgb <= "101111";
					when "010100110000101" => rgb <= "101111";
					when "010100110000110" => rgb <= "101111";
					when "010100110000111" => rgb <= "101111";
					when "010100110001000" => rgb <= "101111";
					when "010100110001001" => rgb <= "101111";
					when "010100110001010" => rgb <= "101111";
					when "010100110001011" => rgb <= "101111";
					when "010100110001100" => rgb <= "101111";
					when "010100110001101" => rgb <= "101111";
					when "010100110001110" => rgb <= "101111";
					when "010100110001111" => rgb <= "101111";
					when "010100110010000" => rgb <= "101111";
					when "010100110010001" => rgb <= "101111";
					when "010100110010010" => rgb <= "101111";
					when "010100110010011" => rgb <= "101111";
					when "010100110010100" => rgb <= "101111";
					when "010100110010101" => rgb <= "101111";
					when "010100110010110" => rgb <= "101111";
					when "010100110010111" => rgb <= "101111";
					when "010100110011000" => rgb <= "101111";
					when "010100110011001" => rgb <= "101111";
					when "010100110011010" => rgb <= "101111";
					when "010100110011011" => rgb <= "101111";
					when "010100110011100" => rgb <= "101111";
					when "010100110011101" => rgb <= "101111";
					when "010100110011110" => rgb <= "101111";
					when "010100110011111" => rgb <= "101111";
					when "010101000000000" => rgb <= "001000";
					when "010101000000001" => rgb <= "001000";
					when "010101000000010" => rgb <= "001000";
					when "010101000000011" => rgb <= "001000";
					when "010101000000100" => rgb <= "001000";
					when "010101000000101" => rgb <= "001000";
					when "010101000000110" => rgb <= "001000";
					when "010101000000111" => rgb <= "001000";
					when "010101000001000" => rgb <= "001000";
					when "010101000001001" => rgb <= "001000";
					when "010101000001010" => rgb <= "001000";
					when "010101000001011" => rgb <= "001000";
					when "010101000001100" => rgb <= "001000";
					when "010101000001101" => rgb <= "001000";
					when "010101000001110" => rgb <= "001000";
					when "010101000001111" => rgb <= "001000";
					when "010101000010000" => rgb <= "001000";
					when "010101000010001" => rgb <= "001000";
					when "010101000010010" => rgb <= "001000";
					when "010101000010011" => rgb <= "001000";
					when "010101000010100" => rgb <= "001000";
					when "010101000010101" => rgb <= "001000";
					when "010101000010110" => rgb <= "001000";
					when "010101000010111" => rgb <= "001000";
					when "010101000011000" => rgb <= "001000";
					when "010101000011001" => rgb <= "001000";
					when "010101000011010" => rgb <= "001000";
					when "010101000011011" => rgb <= "001000";
					when "010101000011100" => rgb <= "001000";
					when "010101000011101" => rgb <= "001000";
					when "010101000011110" => rgb <= "001000";
					when "010101000011111" => rgb <= "001000";
					when "010101000100000" => rgb <= "001000";
					when "010101000100001" => rgb <= "001000";
					when "010101000100010" => rgb <= "001000";
					when "010101000100011" => rgb <= "001000";
					when "010101000100100" => rgb <= "001000";
					when "010101000100101" => rgb <= "001000";
					when "010101000100110" => rgb <= "001000";
					when "010101000100111" => rgb <= "001000";
					when "010101000101000" => rgb <= "001000";
					when "010101000101001" => rgb <= "001000";
					when "010101000101010" => rgb <= "001000";
					when "010101000101011" => rgb <= "001000";
					when "010101000101100" => rgb <= "001000";
					when "010101000101101" => rgb <= "001000";
					when "010101000101110" => rgb <= "001000";
					when "010101000101111" => rgb <= "001000";
					when "010101000110000" => rgb <= "001000";
					when "010101000110001" => rgb <= "001000";
					when "010101000110010" => rgb <= "001000";
					when "010101000110011" => rgb <= "001000";
					when "010101000110100" => rgb <= "001000";
					when "010101000110101" => rgb <= "001000";
					when "010101000110110" => rgb <= "001000";
					when "010101000110111" => rgb <= "001000";
					when "010101000111000" => rgb <= "001000";
					when "010101000111001" => rgb <= "001000";
					when "010101000111010" => rgb <= "001000";
					when "010101000111011" => rgb <= "001000";
					when "010101000111100" => rgb <= "001000";
					when "010101000111101" => rgb <= "001000";
					when "010101000111110" => rgb <= "001000";
					when "010101000111111" => rgb <= "001000";
					when "010101001000000" => rgb <= "001000";
					when "010101001000001" => rgb <= "001000";
					when "010101001000010" => rgb <= "001000";
					when "010101001000011" => rgb <= "001000";
					when "010101001000100" => rgb <= "001000";
					when "010101001000101" => rgb <= "001000";
					when "010101001000110" => rgb <= "001000";
					when "010101001000111" => rgb <= "001000";
					when "010101001001000" => rgb <= "001000";
					when "010101001001001" => rgb <= "001000";
					when "010101001001010" => rgb <= "001000";
					when "010101001001011" => rgb <= "001000";
					when "010101001001100" => rgb <= "001000";
					when "010101001001101" => rgb <= "001000";
					when "010101001001110" => rgb <= "001000";
					when "010101001001111" => rgb <= "001000";
					when "010101001010000" => rgb <= "001000";
					when "010101001010001" => rgb <= "001000";
					when "010101001010010" => rgb <= "001000";
					when "010101001010011" => rgb <= "001000";
					when "010101001010100" => rgb <= "001000";
					when "010101001010101" => rgb <= "001000";
					when "010101001010110" => rgb <= "001000";
					when "010101001010111" => rgb <= "001000";
					when "010101001011000" => rgb <= "000000";
					when "010101001011001" => rgb <= "000000";
					when "010101001011010" => rgb <= "101111";
					when "010101001011011" => rgb <= "101111";
					when "010101001011100" => rgb <= "101111";
					when "010101001011101" => rgb <= "101111";
					when "010101001011110" => rgb <= "101111";
					when "010101001011111" => rgb <= "101111";
					when "010101001100000" => rgb <= "101111";
					when "010101001100001" => rgb <= "101111";
					when "010101001100010" => rgb <= "101111";
					when "010101001100011" => rgb <= "101111";
					when "010101001100100" => rgb <= "101111";
					when "010101001100101" => rgb <= "101111";
					when "010101001100110" => rgb <= "101111";
					when "010101001100111" => rgb <= "101111";
					when "010101001101000" => rgb <= "101111";
					when "010101001101001" => rgb <= "101111";
					when "010101001101010" => rgb <= "101111";
					when "010101001101011" => rgb <= "101111";
					when "010101001101100" => rgb <= "101111";
					when "010101001101101" => rgb <= "101111";
					when "010101001101110" => rgb <= "101111";
					when "010101001101111" => rgb <= "101111";
					when "010101001110000" => rgb <= "101111";
					when "010101001110001" => rgb <= "101111";
					when "010101001110010" => rgb <= "101111";
					when "010101001110011" => rgb <= "101111";
					when "010101001110100" => rgb <= "101111";
					when "010101001110101" => rgb <= "101111";
					when "010101001110110" => rgb <= "101111";
					when "010101001110111" => rgb <= "101111";
					when "010101001111000" => rgb <= "101111";
					when "010101001111001" => rgb <= "101111";
					when "010101001111010" => rgb <= "101111";
					when "010101001111011" => rgb <= "101111";
					when "010101001111100" => rgb <= "101111";
					when "010101001111101" => rgb <= "101111";
					when "010101001111110" => rgb <= "101111";
					when "010101001111111" => rgb <= "101111";
					when "010101010000000" => rgb <= "101111";
					when "010101010000001" => rgb <= "101111";
					when "010101010000010" => rgb <= "101111";
					when "010101010000011" => rgb <= "101111";
					when "010101010000100" => rgb <= "101111";
					when "010101010000101" => rgb <= "101111";
					when "010101010000110" => rgb <= "101111";
					when "010101010000111" => rgb <= "101111";
					when "010101010001000" => rgb <= "101111";
					when "010101010001001" => rgb <= "101111";
					when "010101010001010" => rgb <= "101111";
					when "010101010001011" => rgb <= "101111";
					when "010101010001100" => rgb <= "101111";
					when "010101010001101" => rgb <= "101111";
					when "010101010001110" => rgb <= "101111";
					when "010101010001111" => rgb <= "101111";
					when "010101010010000" => rgb <= "101111";
					when "010101010010001" => rgb <= "101111";
					when "010101010010010" => rgb <= "101111";
					when "010101010010011" => rgb <= "101111";
					when "010101010010100" => rgb <= "101111";
					when "010101010010101" => rgb <= "101111";
					when "010101010010110" => rgb <= "101111";
					when "010101010010111" => rgb <= "101111";
					when "010101010011000" => rgb <= "101111";
					when "010101010011001" => rgb <= "101111";
					when "010101010011010" => rgb <= "101111";
					when "010101010011011" => rgb <= "101111";
					when "010101010011100" => rgb <= "101111";
					when "010101010011101" => rgb <= "101111";
					when "010101010011110" => rgb <= "101111";
					when "010101010011111" => rgb <= "101111";
					when "010101100000000" => rgb <= "001000";
					when "010101100000001" => rgb <= "001000";
					when "010101100000010" => rgb <= "001000";
					when "010101100000011" => rgb <= "001000";
					when "010101100000100" => rgb <= "001000";
					when "010101100000101" => rgb <= "001000";
					when "010101100000110" => rgb <= "001000";
					when "010101100000111" => rgb <= "001000";
					when "010101100001000" => rgb <= "001000";
					when "010101100001001" => rgb <= "001000";
					when "010101100001010" => rgb <= "001000";
					when "010101100001011" => rgb <= "001000";
					when "010101100001100" => rgb <= "001000";
					when "010101100001101" => rgb <= "001000";
					when "010101100001110" => rgb <= "001000";
					when "010101100001111" => rgb <= "001000";
					when "010101100010000" => rgb <= "001000";
					when "010101100010001" => rgb <= "001000";
					when "010101100010010" => rgb <= "001000";
					when "010101100010011" => rgb <= "001000";
					when "010101100010100" => rgb <= "001000";
					when "010101100010101" => rgb <= "001000";
					when "010101100010110" => rgb <= "001000";
					when "010101100010111" => rgb <= "001000";
					when "010101100011000" => rgb <= "001000";
					when "010101100011001" => rgb <= "001000";
					when "010101100011010" => rgb <= "001000";
					when "010101100011011" => rgb <= "001000";
					when "010101100011100" => rgb <= "001000";
					when "010101100011101" => rgb <= "001000";
					when "010101100011110" => rgb <= "001000";
					when "010101100011111" => rgb <= "001000";
					when "010101100100000" => rgb <= "001000";
					when "010101100100001" => rgb <= "001000";
					when "010101100100010" => rgb <= "001000";
					when "010101100100011" => rgb <= "001000";
					when "010101100100100" => rgb <= "001000";
					when "010101100100101" => rgb <= "001000";
					when "010101100100110" => rgb <= "001000";
					when "010101100100111" => rgb <= "001000";
					when "010101100101000" => rgb <= "001000";
					when "010101100101001" => rgb <= "001000";
					when "010101100101010" => rgb <= "001000";
					when "010101100101011" => rgb <= "001000";
					when "010101100101100" => rgb <= "001000";
					when "010101100101101" => rgb <= "001000";
					when "010101100101110" => rgb <= "001000";
					when "010101100101111" => rgb <= "001000";
					when "010101100110000" => rgb <= "001000";
					when "010101100110001" => rgb <= "001000";
					when "010101100110010" => rgb <= "001000";
					when "010101100110011" => rgb <= "001000";
					when "010101100110100" => rgb <= "001000";
					when "010101100110101" => rgb <= "001000";
					when "010101100110110" => rgb <= "001000";
					when "010101100110111" => rgb <= "001000";
					when "010101100111000" => rgb <= "001000";
					when "010101100111001" => rgb <= "001000";
					when "010101100111010" => rgb <= "001000";
					when "010101100111011" => rgb <= "001000";
					when "010101100111100" => rgb <= "001000";
					when "010101100111101" => rgb <= "001000";
					when "010101100111110" => rgb <= "001000";
					when "010101100111111" => rgb <= "001000";
					when "010101101000000" => rgb <= "001000";
					when "010101101000001" => rgb <= "001000";
					when "010101101000010" => rgb <= "001000";
					when "010101101000011" => rgb <= "001000";
					when "010101101000100" => rgb <= "001000";
					when "010101101000101" => rgb <= "001000";
					when "010101101000110" => rgb <= "001000";
					when "010101101000111" => rgb <= "001000";
					when "010101101001000" => rgb <= "001000";
					when "010101101001001" => rgb <= "001000";
					when "010101101001010" => rgb <= "001000";
					when "010101101001011" => rgb <= "001000";
					when "010101101001100" => rgb <= "001000";
					when "010101101001101" => rgb <= "001000";
					when "010101101001110" => rgb <= "001000";
					when "010101101001111" => rgb <= "001000";
					when "010101101010000" => rgb <= "001000";
					when "010101101010001" => rgb <= "001000";
					when "010101101010010" => rgb <= "001000";
					when "010101101010011" => rgb <= "001000";
					when "010101101010100" => rgb <= "001000";
					when "010101101010101" => rgb <= "001000";
					when "010101101010110" => rgb <= "001000";
					when "010101101010111" => rgb <= "001000";
					when "010101101011000" => rgb <= "000000";
					when "010101101011001" => rgb <= "000000";
					when "010101101011010" => rgb <= "101111";
					when "010101101011011" => rgb <= "101111";
					when "010101101011100" => rgb <= "101111";
					when "010101101011101" => rgb <= "101111";
					when "010101101011110" => rgb <= "101111";
					when "010101101011111" => rgb <= "101111";
					when "010101101100000" => rgb <= "101111";
					when "010101101100001" => rgb <= "101111";
					when "010101101100010" => rgb <= "101111";
					when "010101101100011" => rgb <= "101111";
					when "010101101100100" => rgb <= "101111";
					when "010101101100101" => rgb <= "101111";
					when "010101101100110" => rgb <= "101111";
					when "010101101100111" => rgb <= "101111";
					when "010101101101000" => rgb <= "101111";
					when "010101101101001" => rgb <= "101111";
					when "010101101101010" => rgb <= "101111";
					when "010101101101011" => rgb <= "101111";
					when "010101101101100" => rgb <= "101111";
					when "010101101101101" => rgb <= "101111";
					when "010101101101110" => rgb <= "101111";
					when "010101101101111" => rgb <= "101111";
					when "010101101110000" => rgb <= "101111";
					when "010101101110001" => rgb <= "101111";
					when "010101101110010" => rgb <= "101111";
					when "010101101110011" => rgb <= "101111";
					when "010101101110100" => rgb <= "101111";
					when "010101101110101" => rgb <= "101111";
					when "010101101110110" => rgb <= "101111";
					when "010101101110111" => rgb <= "101111";
					when "010101101111000" => rgb <= "101111";
					when "010101101111001" => rgb <= "101111";
					when "010101101111010" => rgb <= "101111";
					when "010101101111011" => rgb <= "101111";
					when "010101101111100" => rgb <= "101111";
					when "010101101111101" => rgb <= "101111";
					when "010101101111110" => rgb <= "101111";
					when "010101101111111" => rgb <= "101111";
					when "010101110000000" => rgb <= "101111";
					when "010101110000001" => rgb <= "101111";
					when "010101110000010" => rgb <= "101111";
					when "010101110000011" => rgb <= "101111";
					when "010101110000100" => rgb <= "101111";
					when "010101110000101" => rgb <= "101111";
					when "010101110000110" => rgb <= "101111";
					when "010101110000111" => rgb <= "101111";
					when "010101110001000" => rgb <= "101111";
					when "010101110001001" => rgb <= "101111";
					when "010101110001010" => rgb <= "101111";
					when "010101110001011" => rgb <= "101111";
					when "010101110001100" => rgb <= "101111";
					when "010101110001101" => rgb <= "101111";
					when "010101110001110" => rgb <= "101111";
					when "010101110001111" => rgb <= "101111";
					when "010101110010000" => rgb <= "101111";
					when "010101110010001" => rgb <= "101111";
					when "010101110010010" => rgb <= "101111";
					when "010101110010011" => rgb <= "101111";
					when "010101110010100" => rgb <= "101111";
					when "010101110010101" => rgb <= "101111";
					when "010101110010110" => rgb <= "101111";
					when "010101110010111" => rgb <= "101111";
					when "010101110011000" => rgb <= "101111";
					when "010101110011001" => rgb <= "101111";
					when "010101110011010" => rgb <= "101111";
					when "010101110011011" => rgb <= "101111";
					when "010101110011100" => rgb <= "101111";
					when "010101110011101" => rgb <= "101111";
					when "010101110011110" => rgb <= "101111";
					when "010101110011111" => rgb <= "101111";
					when "010110000000000" => rgb <= "001000";
					when "010110000000001" => rgb <= "001000";
					when "010110000000010" => rgb <= "001000";
					when "010110000000011" => rgb <= "001000";
					when "010110000000100" => rgb <= "001000";
					when "010110000000101" => rgb <= "001000";
					when "010110000000110" => rgb <= "001000";
					when "010110000000111" => rgb <= "001000";
					when "010110000001000" => rgb <= "001000";
					when "010110000001001" => rgb <= "001000";
					when "010110000001010" => rgb <= "001000";
					when "010110000001011" => rgb <= "001000";
					when "010110000001100" => rgb <= "001000";
					when "010110000001101" => rgb <= "001000";
					when "010110000001110" => rgb <= "001000";
					when "010110000001111" => rgb <= "001000";
					when "010110000010000" => rgb <= "001000";
					when "010110000010001" => rgb <= "001000";
					when "010110000010010" => rgb <= "001000";
					when "010110000010011" => rgb <= "001000";
					when "010110000010100" => rgb <= "001000";
					when "010110000010101" => rgb <= "001000";
					when "010110000010110" => rgb <= "001000";
					when "010110000010111" => rgb <= "001000";
					when "010110000011000" => rgb <= "001000";
					when "010110000011001" => rgb <= "001000";
					when "010110000011010" => rgb <= "001000";
					when "010110000011011" => rgb <= "001000";
					when "010110000011100" => rgb <= "001000";
					when "010110000011101" => rgb <= "001000";
					when "010110000011110" => rgb <= "001000";
					when "010110000011111" => rgb <= "001000";
					when "010110000100000" => rgb <= "001000";
					when "010110000100001" => rgb <= "001000";
					when "010110000100010" => rgb <= "001000";
					when "010110000100011" => rgb <= "001000";
					when "010110000100100" => rgb <= "001000";
					when "010110000100101" => rgb <= "001000";
					when "010110000100110" => rgb <= "001000";
					when "010110000100111" => rgb <= "001000";
					when "010110000101000" => rgb <= "001000";
					when "010110000101001" => rgb <= "001000";
					when "010110000101010" => rgb <= "001000";
					when "010110000101011" => rgb <= "001000";
					when "010110000101100" => rgb <= "001000";
					when "010110000101101" => rgb <= "001000";
					when "010110000101110" => rgb <= "001000";
					when "010110000101111" => rgb <= "001000";
					when "010110000110000" => rgb <= "001000";
					when "010110000110001" => rgb <= "001000";
					when "010110000110010" => rgb <= "001000";
					when "010110000110011" => rgb <= "001000";
					when "010110000110100" => rgb <= "001000";
					when "010110000110101" => rgb <= "001000";
					when "010110000110110" => rgb <= "001000";
					when "010110000110111" => rgb <= "001000";
					when "010110000111000" => rgb <= "001000";
					when "010110000111001" => rgb <= "001000";
					when "010110000111010" => rgb <= "001000";
					when "010110000111011" => rgb <= "001000";
					when "010110000111100" => rgb <= "001000";
					when "010110000111101" => rgb <= "001000";
					when "010110000111110" => rgb <= "001000";
					when "010110000111111" => rgb <= "001000";
					when "010110001000000" => rgb <= "001000";
					when "010110001000001" => rgb <= "001000";
					when "010110001000010" => rgb <= "001000";
					when "010110001000011" => rgb <= "001000";
					when "010110001000100" => rgb <= "001000";
					when "010110001000101" => rgb <= "001000";
					when "010110001000110" => rgb <= "001000";
					when "010110001000111" => rgb <= "001000";
					when "010110001001000" => rgb <= "001000";
					when "010110001001001" => rgb <= "001000";
					when "010110001001010" => rgb <= "001000";
					when "010110001001011" => rgb <= "001000";
					when "010110001001100" => rgb <= "001000";
					when "010110001001101" => rgb <= "001000";
					when "010110001001110" => rgb <= "001000";
					when "010110001001111" => rgb <= "001000";
					when "010110001010000" => rgb <= "001000";
					when "010110001010001" => rgb <= "001000";
					when "010110001010010" => rgb <= "001000";
					when "010110001010011" => rgb <= "001000";
					when "010110001010100" => rgb <= "001000";
					when "010110001010101" => rgb <= "001000";
					when "010110001010110" => rgb <= "000000";
					when "010110001010111" => rgb <= "000000";
					when "010110001011000" => rgb <= "000000";
					when "010110001011001" => rgb <= "000000";
					when "010110001011010" => rgb <= "101111";
					when "010110001011011" => rgb <= "101111";
					when "010110001011100" => rgb <= "101111";
					when "010110001011101" => rgb <= "101111";
					when "010110001011110" => rgb <= "101111";
					when "010110001011111" => rgb <= "101111";
					when "010110001100000" => rgb <= "101111";
					when "010110001100001" => rgb <= "101111";
					when "010110001100010" => rgb <= "101111";
					when "010110001100011" => rgb <= "101111";
					when "010110001100100" => rgb <= "101111";
					when "010110001100101" => rgb <= "101111";
					when "010110001100110" => rgb <= "101111";
					when "010110001100111" => rgb <= "101111";
					when "010110001101000" => rgb <= "101111";
					when "010110001101001" => rgb <= "101111";
					when "010110001101010" => rgb <= "101111";
					when "010110001101011" => rgb <= "101111";
					when "010110001101100" => rgb <= "101111";
					when "010110001101101" => rgb <= "101111";
					when "010110001101110" => rgb <= "101111";
					when "010110001101111" => rgb <= "101111";
					when "010110001110000" => rgb <= "101111";
					when "010110001110001" => rgb <= "101111";
					when "010110001110010" => rgb <= "101111";
					when "010110001110011" => rgb <= "101111";
					when "010110001110100" => rgb <= "101111";
					when "010110001110101" => rgb <= "101111";
					when "010110001110110" => rgb <= "101111";
					when "010110001110111" => rgb <= "101111";
					when "010110001111000" => rgb <= "101111";
					when "010110001111001" => rgb <= "101111";
					when "010110001111010" => rgb <= "101111";
					when "010110001111011" => rgb <= "101111";
					when "010110001111100" => rgb <= "101111";
					when "010110001111101" => rgb <= "101111";
					when "010110001111110" => rgb <= "101111";
					when "010110001111111" => rgb <= "101111";
					when "010110010000000" => rgb <= "101111";
					when "010110010000001" => rgb <= "101111";
					when "010110010000010" => rgb <= "101111";
					when "010110010000011" => rgb <= "101111";
					when "010110010000100" => rgb <= "101111";
					when "010110010000101" => rgb <= "101111";
					when "010110010000110" => rgb <= "101111";
					when "010110010000111" => rgb <= "101111";
					when "010110010001000" => rgb <= "101111";
					when "010110010001001" => rgb <= "101111";
					when "010110010001010" => rgb <= "101111";
					when "010110010001011" => rgb <= "101111";
					when "010110010001100" => rgb <= "101111";
					when "010110010001101" => rgb <= "101111";
					when "010110010001110" => rgb <= "101111";
					when "010110010001111" => rgb <= "101111";
					when "010110010010000" => rgb <= "101111";
					when "010110010010001" => rgb <= "101111";
					when "010110010010010" => rgb <= "101111";
					when "010110010010011" => rgb <= "101111";
					when "010110010010100" => rgb <= "101111";
					when "010110010010101" => rgb <= "101111";
					when "010110010010110" => rgb <= "101111";
					when "010110010010111" => rgb <= "101111";
					when "010110010011000" => rgb <= "101111";
					when "010110010011001" => rgb <= "101111";
					when "010110010011010" => rgb <= "101111";
					when "010110010011011" => rgb <= "101111";
					when "010110010011100" => rgb <= "101111";
					when "010110010011101" => rgb <= "101111";
					when "010110010011110" => rgb <= "101111";
					when "010110010011111" => rgb <= "101111";
					when "010110100000000" => rgb <= "001000";
					when "010110100000001" => rgb <= "001000";
					when "010110100000010" => rgb <= "001000";
					when "010110100000011" => rgb <= "001000";
					when "010110100000100" => rgb <= "001000";
					when "010110100000101" => rgb <= "001000";
					when "010110100000110" => rgb <= "001000";
					when "010110100000111" => rgb <= "001000";
					when "010110100001000" => rgb <= "001000";
					when "010110100001001" => rgb <= "001000";
					when "010110100001010" => rgb <= "001000";
					when "010110100001011" => rgb <= "001000";
					when "010110100001100" => rgb <= "001000";
					when "010110100001101" => rgb <= "001000";
					when "010110100001110" => rgb <= "001000";
					when "010110100001111" => rgb <= "001000";
					when "010110100010000" => rgb <= "001000";
					when "010110100010001" => rgb <= "001000";
					when "010110100010010" => rgb <= "001000";
					when "010110100010011" => rgb <= "001000";
					when "010110100010100" => rgb <= "001000";
					when "010110100010101" => rgb <= "001000";
					when "010110100010110" => rgb <= "001000";
					when "010110100010111" => rgb <= "001000";
					when "010110100011000" => rgb <= "001000";
					when "010110100011001" => rgb <= "001000";
					when "010110100011010" => rgb <= "001000";
					when "010110100011011" => rgb <= "001000";
					when "010110100011100" => rgb <= "001000";
					when "010110100011101" => rgb <= "001000";
					when "010110100011110" => rgb <= "001000";
					when "010110100011111" => rgb <= "001000";
					when "010110100100000" => rgb <= "001000";
					when "010110100100001" => rgb <= "001000";
					when "010110100100010" => rgb <= "001000";
					when "010110100100011" => rgb <= "001000";
					when "010110100100100" => rgb <= "001000";
					when "010110100100101" => rgb <= "001000";
					when "010110100100110" => rgb <= "001000";
					when "010110100100111" => rgb <= "001000";
					when "010110100101000" => rgb <= "001000";
					when "010110100101001" => rgb <= "001000";
					when "010110100101010" => rgb <= "001000";
					when "010110100101011" => rgb <= "001000";
					when "010110100101100" => rgb <= "001000";
					when "010110100101101" => rgb <= "001000";
					when "010110100101110" => rgb <= "001000";
					when "010110100101111" => rgb <= "001000";
					when "010110100110000" => rgb <= "001000";
					when "010110100110001" => rgb <= "001000";
					when "010110100110010" => rgb <= "001000";
					when "010110100110011" => rgb <= "001000";
					when "010110100110100" => rgb <= "001000";
					when "010110100110101" => rgb <= "001000";
					when "010110100110110" => rgb <= "001000";
					when "010110100110111" => rgb <= "001000";
					when "010110100111000" => rgb <= "001000";
					when "010110100111001" => rgb <= "001000";
					when "010110100111010" => rgb <= "001000";
					when "010110100111011" => rgb <= "001000";
					when "010110100111100" => rgb <= "001000";
					when "010110100111101" => rgb <= "001000";
					when "010110100111110" => rgb <= "001000";
					when "010110100111111" => rgb <= "001000";
					when "010110101000000" => rgb <= "001000";
					when "010110101000001" => rgb <= "001000";
					when "010110101000010" => rgb <= "001000";
					when "010110101000011" => rgb <= "001000";
					when "010110101000100" => rgb <= "001000";
					when "010110101000101" => rgb <= "001000";
					when "010110101000110" => rgb <= "001000";
					when "010110101000111" => rgb <= "001000";
					when "010110101001000" => rgb <= "001000";
					when "010110101001001" => rgb <= "001000";
					when "010110101001010" => rgb <= "001000";
					when "010110101001011" => rgb <= "001000";
					when "010110101001100" => rgb <= "001000";
					when "010110101001101" => rgb <= "001000";
					when "010110101001110" => rgb <= "001000";
					when "010110101001111" => rgb <= "001000";
					when "010110101010000" => rgb <= "001000";
					when "010110101010001" => rgb <= "001000";
					when "010110101010010" => rgb <= "001000";
					when "010110101010011" => rgb <= "001000";
					when "010110101010100" => rgb <= "001000";
					when "010110101010101" => rgb <= "001000";
					when "010110101010110" => rgb <= "000000";
					when "010110101010111" => rgb <= "000000";
					when "010110101011000" => rgb <= "000000";
					when "010110101011001" => rgb <= "000000";
					when "010110101011010" => rgb <= "101111";
					when "010110101011011" => rgb <= "101111";
					when "010110101011100" => rgb <= "101111";
					when "010110101011101" => rgb <= "101111";
					when "010110101011110" => rgb <= "101111";
					when "010110101011111" => rgb <= "101111";
					when "010110101100000" => rgb <= "101111";
					when "010110101100001" => rgb <= "101111";
					when "010110101100010" => rgb <= "101111";
					when "010110101100011" => rgb <= "101111";
					when "010110101100100" => rgb <= "101111";
					when "010110101100101" => rgb <= "101111";
					when "010110101100110" => rgb <= "101111";
					when "010110101100111" => rgb <= "101111";
					when "010110101101000" => rgb <= "101111";
					when "010110101101001" => rgb <= "101111";
					when "010110101101010" => rgb <= "101111";
					when "010110101101011" => rgb <= "101111";
					when "010110101101100" => rgb <= "101111";
					when "010110101101101" => rgb <= "101111";
					when "010110101101110" => rgb <= "101111";
					when "010110101101111" => rgb <= "101111";
					when "010110101110000" => rgb <= "101111";
					when "010110101110001" => rgb <= "101111";
					when "010110101110010" => rgb <= "101111";
					when "010110101110011" => rgb <= "101111";
					when "010110101110100" => rgb <= "101111";
					when "010110101110101" => rgb <= "101111";
					when "010110101110110" => rgb <= "101111";
					when "010110101110111" => rgb <= "101111";
					when "010110101111000" => rgb <= "101111";
					when "010110101111001" => rgb <= "101111";
					when "010110101111010" => rgb <= "101111";
					when "010110101111011" => rgb <= "101111";
					when "010110101111100" => rgb <= "101111";
					when "010110101111101" => rgb <= "101111";
					when "010110101111110" => rgb <= "101111";
					when "010110101111111" => rgb <= "101111";
					when "010110110000000" => rgb <= "101111";
					when "010110110000001" => rgb <= "101111";
					when "010110110000010" => rgb <= "101111";
					when "010110110000011" => rgb <= "101111";
					when "010110110000100" => rgb <= "101111";
					when "010110110000101" => rgb <= "101111";
					when "010110110000110" => rgb <= "101111";
					when "010110110000111" => rgb <= "101111";
					when "010110110001000" => rgb <= "101111";
					when "010110110001001" => rgb <= "101111";
					when "010110110001010" => rgb <= "101111";
					when "010110110001011" => rgb <= "101111";
					when "010110110001100" => rgb <= "101111";
					when "010110110001101" => rgb <= "101111";
					when "010110110001110" => rgb <= "101111";
					when "010110110001111" => rgb <= "101111";
					when "010110110010000" => rgb <= "101111";
					when "010110110010001" => rgb <= "101111";
					when "010110110010010" => rgb <= "101111";
					when "010110110010011" => rgb <= "101111";
					when "010110110010100" => rgb <= "101111";
					when "010110110010101" => rgb <= "101111";
					when "010110110010110" => rgb <= "101111";
					when "010110110010111" => rgb <= "101111";
					when "010110110011000" => rgb <= "101111";
					when "010110110011001" => rgb <= "101111";
					when "010110110011010" => rgb <= "101111";
					when "010110110011011" => rgb <= "101111";
					when "010110110011100" => rgb <= "101111";
					when "010110110011101" => rgb <= "101111";
					when "010110110011110" => rgb <= "101111";
					when "010110110011111" => rgb <= "101111";
					when "010111000000000" => rgb <= "001000";
					when "010111000000001" => rgb <= "001000";
					when "010111000000010" => rgb <= "001000";
					when "010111000000011" => rgb <= "001000";
					when "010111000000100" => rgb <= "001000";
					when "010111000000101" => rgb <= "001000";
					when "010111000000110" => rgb <= "001000";
					when "010111000000111" => rgb <= "001000";
					when "010111000001000" => rgb <= "001000";
					when "010111000001001" => rgb <= "001000";
					when "010111000001010" => rgb <= "001000";
					when "010111000001011" => rgb <= "001000";
					when "010111000001100" => rgb <= "001000";
					when "010111000001101" => rgb <= "001000";
					when "010111000001110" => rgb <= "001000";
					when "010111000001111" => rgb <= "001000";
					when "010111000010000" => rgb <= "001000";
					when "010111000010001" => rgb <= "001000";
					when "010111000010010" => rgb <= "001000";
					when "010111000010011" => rgb <= "001000";
					when "010111000010100" => rgb <= "001000";
					when "010111000010101" => rgb <= "001000";
					when "010111000010110" => rgb <= "001000";
					when "010111000010111" => rgb <= "001000";
					when "010111000011000" => rgb <= "001000";
					when "010111000011001" => rgb <= "001000";
					when "010111000011010" => rgb <= "001000";
					when "010111000011011" => rgb <= "001000";
					when "010111000011100" => rgb <= "001000";
					when "010111000011101" => rgb <= "001000";
					when "010111000011110" => rgb <= "001000";
					when "010111000011111" => rgb <= "001000";
					when "010111000100000" => rgb <= "001000";
					when "010111000100001" => rgb <= "001000";
					when "010111000100010" => rgb <= "001000";
					when "010111000100011" => rgb <= "001000";
					when "010111000100100" => rgb <= "001000";
					when "010111000100101" => rgb <= "001000";
					when "010111000100110" => rgb <= "001000";
					when "010111000100111" => rgb <= "001000";
					when "010111000101000" => rgb <= "001000";
					when "010111000101001" => rgb <= "001000";
					when "010111000101010" => rgb <= "001000";
					when "010111000101011" => rgb <= "001000";
					when "010111000101100" => rgb <= "001000";
					when "010111000101101" => rgb <= "001000";
					when "010111000101110" => rgb <= "001000";
					when "010111000101111" => rgb <= "001000";
					when "010111000110000" => rgb <= "001000";
					when "010111000110001" => rgb <= "001000";
					when "010111000110010" => rgb <= "001000";
					when "010111000110011" => rgb <= "001000";
					when "010111000110100" => rgb <= "001000";
					when "010111000110101" => rgb <= "001000";
					when "010111000110110" => rgb <= "001000";
					when "010111000110111" => rgb <= "001000";
					when "010111000111000" => rgb <= "001000";
					when "010111000111001" => rgb <= "001000";
					when "010111000111010" => rgb <= "001000";
					when "010111000111011" => rgb <= "001000";
					when "010111000111100" => rgb <= "001000";
					when "010111000111101" => rgb <= "001000";
					when "010111000111110" => rgb <= "001000";
					when "010111000111111" => rgb <= "001000";
					when "010111001000000" => rgb <= "001000";
					when "010111001000001" => rgb <= "001000";
					when "010111001000010" => rgb <= "001000";
					when "010111001000011" => rgb <= "001000";
					when "010111001000100" => rgb <= "001000";
					when "010111001000101" => rgb <= "001000";
					when "010111001000110" => rgb <= "001000";
					when "010111001000111" => rgb <= "001000";
					when "010111001001000" => rgb <= "001000";
					when "010111001001001" => rgb <= "001000";
					when "010111001001010" => rgb <= "001000";
					when "010111001001011" => rgb <= "001000";
					when "010111001001100" => rgb <= "001000";
					when "010111001001101" => rgb <= "001000";
					when "010111001001110" => rgb <= "001000";
					when "010111001001111" => rgb <= "001000";
					when "010111001010000" => rgb <= "001000";
					when "010111001010001" => rgb <= "001000";
					when "010111001010010" => rgb <= "001000";
					when "010111001010011" => rgb <= "001000";
					when "010111001010100" => rgb <= "000000";
					when "010111001010101" => rgb <= "000000";
					when "010111001010110" => rgb <= "101111";
					when "010111001010111" => rgb <= "101111";
					when "010111001011000" => rgb <= "101111";
					when "010111001011001" => rgb <= "101111";
					when "010111001011010" => rgb <= "101111";
					when "010111001011011" => rgb <= "101111";
					when "010111001011100" => rgb <= "101111";
					when "010111001011101" => rgb <= "101111";
					when "010111001011110" => rgb <= "101111";
					when "010111001011111" => rgb <= "101111";
					when "010111001100000" => rgb <= "101111";
					when "010111001100001" => rgb <= "101111";
					when "010111001100010" => rgb <= "101111";
					when "010111001100011" => rgb <= "101111";
					when "010111001100100" => rgb <= "101111";
					when "010111001100101" => rgb <= "101111";
					when "010111001100110" => rgb <= "101111";
					when "010111001100111" => rgb <= "101111";
					when "010111001101000" => rgb <= "101111";
					when "010111001101001" => rgb <= "101111";
					when "010111001101010" => rgb <= "101111";
					when "010111001101011" => rgb <= "101111";
					when "010111001101100" => rgb <= "101111";
					when "010111001101101" => rgb <= "101111";
					when "010111001101110" => rgb <= "101111";
					when "010111001101111" => rgb <= "101111";
					when "010111001110000" => rgb <= "101111";
					when "010111001110001" => rgb <= "101111";
					when "010111001110010" => rgb <= "101111";
					when "010111001110011" => rgb <= "101111";
					when "010111001110100" => rgb <= "101111";
					when "010111001110101" => rgb <= "101111";
					when "010111001110110" => rgb <= "101111";
					when "010111001110111" => rgb <= "101111";
					when "010111001111000" => rgb <= "101111";
					when "010111001111001" => rgb <= "101111";
					when "010111001111010" => rgb <= "101111";
					when "010111001111011" => rgb <= "101111";
					when "010111001111100" => rgb <= "101111";
					when "010111001111101" => rgb <= "101111";
					when "010111001111110" => rgb <= "101111";
					when "010111001111111" => rgb <= "101111";
					when "010111010000000" => rgb <= "101111";
					when "010111010000001" => rgb <= "101111";
					when "010111010000010" => rgb <= "101111";
					when "010111010000011" => rgb <= "101111";
					when "010111010000100" => rgb <= "101111";
					when "010111010000101" => rgb <= "101111";
					when "010111010000110" => rgb <= "101111";
					when "010111010000111" => rgb <= "101111";
					when "010111010001000" => rgb <= "101111";
					when "010111010001001" => rgb <= "101111";
					when "010111010001010" => rgb <= "101111";
					when "010111010001011" => rgb <= "101111";
					when "010111010001100" => rgb <= "101111";
					when "010111010001101" => rgb <= "101111";
					when "010111010001110" => rgb <= "101111";
					when "010111010001111" => rgb <= "101111";
					when "010111010010000" => rgb <= "101111";
					when "010111010010001" => rgb <= "101111";
					when "010111010010010" => rgb <= "101111";
					when "010111010010011" => rgb <= "101111";
					when "010111010010100" => rgb <= "101111";
					when "010111010010101" => rgb <= "101111";
					when "010111010010110" => rgb <= "101111";
					when "010111010010111" => rgb <= "101111";
					when "010111010011000" => rgb <= "101111";
					when "010111010011001" => rgb <= "101111";
					when "010111010011010" => rgb <= "101111";
					when "010111010011011" => rgb <= "101111";
					when "010111010011100" => rgb <= "101111";
					when "010111010011101" => rgb <= "101111";
					when "010111010011110" => rgb <= "101111";
					when "010111010011111" => rgb <= "101111";
					when "010111100000000" => rgb <= "001000";
					when "010111100000001" => rgb <= "001000";
					when "010111100000010" => rgb <= "001000";
					when "010111100000011" => rgb <= "001000";
					when "010111100000100" => rgb <= "001000";
					when "010111100000101" => rgb <= "001000";
					when "010111100000110" => rgb <= "001000";
					when "010111100000111" => rgb <= "001000";
					when "010111100001000" => rgb <= "001000";
					when "010111100001001" => rgb <= "001000";
					when "010111100001010" => rgb <= "001000";
					when "010111100001011" => rgb <= "001000";
					when "010111100001100" => rgb <= "001000";
					when "010111100001101" => rgb <= "001000";
					when "010111100001110" => rgb <= "001000";
					when "010111100001111" => rgb <= "001000";
					when "010111100010000" => rgb <= "001000";
					when "010111100010001" => rgb <= "001000";
					when "010111100010010" => rgb <= "001000";
					when "010111100010011" => rgb <= "001000";
					when "010111100010100" => rgb <= "001000";
					when "010111100010101" => rgb <= "001000";
					when "010111100010110" => rgb <= "001000";
					when "010111100010111" => rgb <= "001000";
					when "010111100011000" => rgb <= "001000";
					when "010111100011001" => rgb <= "001000";
					when "010111100011010" => rgb <= "001000";
					when "010111100011011" => rgb <= "001000";
					when "010111100011100" => rgb <= "001000";
					when "010111100011101" => rgb <= "001000";
					when "010111100011110" => rgb <= "001000";
					when "010111100011111" => rgb <= "001000";
					when "010111100100000" => rgb <= "001000";
					when "010111100100001" => rgb <= "001000";
					when "010111100100010" => rgb <= "001000";
					when "010111100100011" => rgb <= "001000";
					when "010111100100100" => rgb <= "001000";
					when "010111100100101" => rgb <= "001000";
					when "010111100100110" => rgb <= "001000";
					when "010111100100111" => rgb <= "001000";
					when "010111100101000" => rgb <= "001000";
					when "010111100101001" => rgb <= "001000";
					when "010111100101010" => rgb <= "001000";
					when "010111100101011" => rgb <= "001000";
					when "010111100101100" => rgb <= "001000";
					when "010111100101101" => rgb <= "001000";
					when "010111100101110" => rgb <= "001000";
					when "010111100101111" => rgb <= "001000";
					when "010111100110000" => rgb <= "001000";
					when "010111100110001" => rgb <= "001000";
					when "010111100110010" => rgb <= "001000";
					when "010111100110011" => rgb <= "001000";
					when "010111100110100" => rgb <= "001000";
					when "010111100110101" => rgb <= "001000";
					when "010111100110110" => rgb <= "001000";
					when "010111100110111" => rgb <= "001000";
					when "010111100111000" => rgb <= "001000";
					when "010111100111001" => rgb <= "001000";
					when "010111100111010" => rgb <= "001000";
					when "010111100111011" => rgb <= "001000";
					when "010111100111100" => rgb <= "001000";
					when "010111100111101" => rgb <= "001000";
					when "010111100111110" => rgb <= "001000";
					when "010111100111111" => rgb <= "001000";
					when "010111101000000" => rgb <= "001000";
					when "010111101000001" => rgb <= "001000";
					when "010111101000010" => rgb <= "001000";
					when "010111101000011" => rgb <= "001000";
					when "010111101000100" => rgb <= "001000";
					when "010111101000101" => rgb <= "001000";
					when "010111101000110" => rgb <= "001000";
					when "010111101000111" => rgb <= "001000";
					when "010111101001000" => rgb <= "001000";
					when "010111101001001" => rgb <= "001000";
					when "010111101001010" => rgb <= "001000";
					when "010111101001011" => rgb <= "001000";
					when "010111101001100" => rgb <= "001000";
					when "010111101001101" => rgb <= "001000";
					when "010111101001110" => rgb <= "001000";
					when "010111101001111" => rgb <= "001000";
					when "010111101010000" => rgb <= "001000";
					when "010111101010001" => rgb <= "001000";
					when "010111101010010" => rgb <= "001000";
					when "010111101010011" => rgb <= "001000";
					when "010111101010100" => rgb <= "000000";
					when "010111101010101" => rgb <= "000000";
					when "010111101010110" => rgb <= "101111";
					when "010111101010111" => rgb <= "101111";
					when "010111101011000" => rgb <= "101111";
					when "010111101011001" => rgb <= "101111";
					when "010111101011010" => rgb <= "101111";
					when "010111101011011" => rgb <= "101111";
					when "010111101011100" => rgb <= "101111";
					when "010111101011101" => rgb <= "101111";
					when "010111101011110" => rgb <= "101111";
					when "010111101011111" => rgb <= "101111";
					when "010111101100000" => rgb <= "101111";
					when "010111101100001" => rgb <= "101111";
					when "010111101100010" => rgb <= "101111";
					when "010111101100011" => rgb <= "101111";
					when "010111101100100" => rgb <= "101111";
					when "010111101100101" => rgb <= "101111";
					when "010111101100110" => rgb <= "101111";
					when "010111101100111" => rgb <= "101111";
					when "010111101101000" => rgb <= "101111";
					when "010111101101001" => rgb <= "101111";
					when "010111101101010" => rgb <= "101111";
					when "010111101101011" => rgb <= "101111";
					when "010111101101100" => rgb <= "101111";
					when "010111101101101" => rgb <= "101111";
					when "010111101101110" => rgb <= "101111";
					when "010111101101111" => rgb <= "101111";
					when "010111101110000" => rgb <= "101111";
					when "010111101110001" => rgb <= "101111";
					when "010111101110010" => rgb <= "101111";
					when "010111101110011" => rgb <= "101111";
					when "010111101110100" => rgb <= "101111";
					when "010111101110101" => rgb <= "101111";
					when "010111101110110" => rgb <= "101111";
					when "010111101110111" => rgb <= "101111";
					when "010111101111000" => rgb <= "101111";
					when "010111101111001" => rgb <= "101111";
					when "010111101111010" => rgb <= "101111";
					when "010111101111011" => rgb <= "101111";
					when "010111101111100" => rgb <= "101111";
					when "010111101111101" => rgb <= "101111";
					when "010111101111110" => rgb <= "101111";
					when "010111101111111" => rgb <= "101111";
					when "010111110000000" => rgb <= "101111";
					when "010111110000001" => rgb <= "101111";
					when "010111110000010" => rgb <= "101111";
					when "010111110000011" => rgb <= "101111";
					when "010111110000100" => rgb <= "101111";
					when "010111110000101" => rgb <= "101111";
					when "010111110000110" => rgb <= "101111";
					when "010111110000111" => rgb <= "101111";
					when "010111110001000" => rgb <= "101111";
					when "010111110001001" => rgb <= "101111";
					when "010111110001010" => rgb <= "101111";
					when "010111110001011" => rgb <= "101111";
					when "010111110001100" => rgb <= "101111";
					when "010111110001101" => rgb <= "101111";
					when "010111110001110" => rgb <= "101111";
					when "010111110001111" => rgb <= "101111";
					when "010111110010000" => rgb <= "101111";
					when "010111110010001" => rgb <= "101111";
					when "010111110010010" => rgb <= "101111";
					when "010111110010011" => rgb <= "101111";
					when "010111110010100" => rgb <= "101111";
					when "010111110010101" => rgb <= "101111";
					when "010111110010110" => rgb <= "101111";
					when "010111110010111" => rgb <= "101111";
					when "010111110011000" => rgb <= "101111";
					when "010111110011001" => rgb <= "101111";
					when "010111110011010" => rgb <= "101111";
					when "010111110011011" => rgb <= "101111";
					when "010111110011100" => rgb <= "101111";
					when "010111110011101" => rgb <= "101111";
					when "010111110011110" => rgb <= "101111";
					when "010111110011111" => rgb <= "101111";
					when "011000000000000" => rgb <= "001000";
					when "011000000000001" => rgb <= "001000";
					when "011000000000010" => rgb <= "001000";
					when "011000000000011" => rgb <= "001000";
					when "011000000000100" => rgb <= "001000";
					when "011000000000101" => rgb <= "001000";
					when "011000000000110" => rgb <= "001000";
					when "011000000000111" => rgb <= "001000";
					when "011000000001000" => rgb <= "001000";
					when "011000000001001" => rgb <= "001000";
					when "011000000001010" => rgb <= "001000";
					when "011000000001011" => rgb <= "001000";
					when "011000000001100" => rgb <= "001000";
					when "011000000001101" => rgb <= "001000";
					when "011000000001110" => rgb <= "001000";
					when "011000000001111" => rgb <= "001000";
					when "011000000010000" => rgb <= "001000";
					when "011000000010001" => rgb <= "001000";
					when "011000000010010" => rgb <= "001000";
					when "011000000010011" => rgb <= "001000";
					when "011000000010100" => rgb <= "001000";
					when "011000000010101" => rgb <= "001000";
					when "011000000010110" => rgb <= "001000";
					when "011000000010111" => rgb <= "001000";
					when "011000000011000" => rgb <= "001000";
					when "011000000011001" => rgb <= "001000";
					when "011000000011010" => rgb <= "001000";
					when "011000000011011" => rgb <= "001000";
					when "011000000011100" => rgb <= "001000";
					when "011000000011101" => rgb <= "001000";
					when "011000000011110" => rgb <= "001000";
					when "011000000011111" => rgb <= "001000";
					when "011000000100000" => rgb <= "001000";
					when "011000000100001" => rgb <= "001000";
					when "011000000100010" => rgb <= "001000";
					when "011000000100011" => rgb <= "001000";
					when "011000000100100" => rgb <= "001000";
					when "011000000100101" => rgb <= "001000";
					when "011000000100110" => rgb <= "001000";
					when "011000000100111" => rgb <= "001000";
					when "011000000101000" => rgb <= "001000";
					when "011000000101001" => rgb <= "001000";
					when "011000000101010" => rgb <= "001000";
					when "011000000101011" => rgb <= "001000";
					when "011000000101100" => rgb <= "001000";
					when "011000000101101" => rgb <= "001000";
					when "011000000101110" => rgb <= "001000";
					when "011000000101111" => rgb <= "001000";
					when "011000000110000" => rgb <= "001000";
					when "011000000110001" => rgb <= "001000";
					when "011000000110010" => rgb <= "001000";
					when "011000000110011" => rgb <= "001000";
					when "011000000110100" => rgb <= "001000";
					when "011000000110101" => rgb <= "001000";
					when "011000000110110" => rgb <= "001000";
					when "011000000110111" => rgb <= "001000";
					when "011000000111000" => rgb <= "001000";
					when "011000000111001" => rgb <= "001000";
					when "011000000111010" => rgb <= "001000";
					when "011000000111011" => rgb <= "001000";
					when "011000000111100" => rgb <= "001000";
					when "011000000111101" => rgb <= "001000";
					when "011000000111110" => rgb <= "001000";
					when "011000000111111" => rgb <= "001000";
					when "011000001000000" => rgb <= "001000";
					when "011000001000001" => rgb <= "001000";
					when "011000001000010" => rgb <= "001000";
					when "011000001000011" => rgb <= "001000";
					when "011000001000100" => rgb <= "001000";
					when "011000001000101" => rgb <= "001000";
					when "011000001000110" => rgb <= "001000";
					when "011000001000111" => rgb <= "001000";
					when "011000001001000" => rgb <= "001000";
					when "011000001001001" => rgb <= "001000";
					when "011000001001010" => rgb <= "001000";
					when "011000001001011" => rgb <= "001000";
					when "011000001001100" => rgb <= "001000";
					when "011000001001101" => rgb <= "001000";
					when "011000001001110" => rgb <= "001000";
					when "011000001001111" => rgb <= "001000";
					when "011000001010000" => rgb <= "001000";
					when "011000001010001" => rgb <= "001000";
					when "011000001010010" => rgb <= "001000";
					when "011000001010011" => rgb <= "001000";
					when "011000001010100" => rgb <= "000000";
					when "011000001010101" => rgb <= "000000";
					when "011000001010110" => rgb <= "101111";
					when "011000001010111" => rgb <= "101111";
					when "011000001011000" => rgb <= "101111";
					when "011000001011001" => rgb <= "101111";
					when "011000001011010" => rgb <= "101111";
					when "011000001011011" => rgb <= "101111";
					when "011000001011100" => rgb <= "101111";
					when "011000001011101" => rgb <= "101111";
					when "011000001011110" => rgb <= "101111";
					when "011000001011111" => rgb <= "101111";
					when "011000001100000" => rgb <= "101111";
					when "011000001100001" => rgb <= "101111";
					when "011000001100010" => rgb <= "101111";
					when "011000001100011" => rgb <= "101111";
					when "011000001100100" => rgb <= "101111";
					when "011000001100101" => rgb <= "101111";
					when "011000001100110" => rgb <= "101111";
					when "011000001100111" => rgb <= "101111";
					when "011000001101000" => rgb <= "101111";
					when "011000001101001" => rgb <= "101111";
					when "011000001101010" => rgb <= "101111";
					when "011000001101011" => rgb <= "101111";
					when "011000001101100" => rgb <= "101111";
					when "011000001101101" => rgb <= "101111";
					when "011000001101110" => rgb <= "101111";
					when "011000001101111" => rgb <= "101111";
					when "011000001110000" => rgb <= "101111";
					when "011000001110001" => rgb <= "101111";
					when "011000001110010" => rgb <= "101111";
					when "011000001110011" => rgb <= "101111";
					when "011000001110100" => rgb <= "101111";
					when "011000001110101" => rgb <= "101111";
					when "011000001110110" => rgb <= "101111";
					when "011000001110111" => rgb <= "101111";
					when "011000001111000" => rgb <= "101111";
					when "011000001111001" => rgb <= "101111";
					when "011000001111010" => rgb <= "101111";
					when "011000001111011" => rgb <= "101111";
					when "011000001111100" => rgb <= "101111";
					when "011000001111101" => rgb <= "101111";
					when "011000001111110" => rgb <= "101111";
					when "011000001111111" => rgb <= "101111";
					when "011000010000000" => rgb <= "101111";
					when "011000010000001" => rgb <= "101111";
					when "011000010000010" => rgb <= "101111";
					when "011000010000011" => rgb <= "101111";
					when "011000010000100" => rgb <= "101111";
					when "011000010000101" => rgb <= "101111";
					when "011000010000110" => rgb <= "101111";
					when "011000010000111" => rgb <= "101111";
					when "011000010001000" => rgb <= "101111";
					when "011000010001001" => rgb <= "101111";
					when "011000010001010" => rgb <= "101111";
					when "011000010001011" => rgb <= "101111";
					when "011000010001100" => rgb <= "101111";
					when "011000010001101" => rgb <= "101111";
					when "011000010001110" => rgb <= "101111";
					when "011000010001111" => rgb <= "101111";
					when "011000010010000" => rgb <= "101111";
					when "011000010010001" => rgb <= "101111";
					when "011000010010010" => rgb <= "101111";
					when "011000010010011" => rgb <= "101111";
					when "011000010010100" => rgb <= "101111";
					when "011000010010101" => rgb <= "101111";
					when "011000010010110" => rgb <= "101111";
					when "011000010010111" => rgb <= "101111";
					when "011000010011000" => rgb <= "101111";
					when "011000010011001" => rgb <= "101111";
					when "011000010011010" => rgb <= "101111";
					when "011000010011011" => rgb <= "101111";
					when "011000010011100" => rgb <= "101111";
					when "011000010011101" => rgb <= "101111";
					when "011000010011110" => rgb <= "101111";
					when "011000010011111" => rgb <= "101111";
					when "011000100000000" => rgb <= "001000";
					when "011000100000001" => rgb <= "001000";
					when "011000100000010" => rgb <= "001000";
					when "011000100000011" => rgb <= "001000";
					when "011000100000100" => rgb <= "001000";
					when "011000100000101" => rgb <= "001000";
					when "011000100000110" => rgb <= "001000";
					when "011000100000111" => rgb <= "001000";
					when "011000100001000" => rgb <= "001000";
					when "011000100001001" => rgb <= "001000";
					when "011000100001010" => rgb <= "001000";
					when "011000100001011" => rgb <= "001000";
					when "011000100001100" => rgb <= "001000";
					when "011000100001101" => rgb <= "001000";
					when "011000100001110" => rgb <= "001000";
					when "011000100001111" => rgb <= "001000";
					when "011000100010000" => rgb <= "001000";
					when "011000100010001" => rgb <= "001000";
					when "011000100010010" => rgb <= "001000";
					when "011000100010011" => rgb <= "001000";
					when "011000100010100" => rgb <= "001000";
					when "011000100010101" => rgb <= "001000";
					when "011000100010110" => rgb <= "001000";
					when "011000100010111" => rgb <= "001000";
					when "011000100011000" => rgb <= "001000";
					when "011000100011001" => rgb <= "001000";
					when "011000100011010" => rgb <= "001000";
					when "011000100011011" => rgb <= "001000";
					when "011000100011100" => rgb <= "001000";
					when "011000100011101" => rgb <= "001000";
					when "011000100011110" => rgb <= "001000";
					when "011000100011111" => rgb <= "001000";
					when "011000100100000" => rgb <= "001000";
					when "011000100100001" => rgb <= "001000";
					when "011000100100010" => rgb <= "001000";
					when "011000100100011" => rgb <= "001000";
					when "011000100100100" => rgb <= "001000";
					when "011000100100101" => rgb <= "001000";
					when "011000100100110" => rgb <= "001000";
					when "011000100100111" => rgb <= "001000";
					when "011000100101000" => rgb <= "001000";
					when "011000100101001" => rgb <= "001000";
					when "011000100101010" => rgb <= "001000";
					when "011000100101011" => rgb <= "001000";
					when "011000100101100" => rgb <= "001000";
					when "011000100101101" => rgb <= "001000";
					when "011000100101110" => rgb <= "001000";
					when "011000100101111" => rgb <= "001000";
					when "011000100110000" => rgb <= "001000";
					when "011000100110001" => rgb <= "001000";
					when "011000100110010" => rgb <= "001000";
					when "011000100110011" => rgb <= "001000";
					when "011000100110100" => rgb <= "001000";
					when "011000100110101" => rgb <= "001000";
					when "011000100110110" => rgb <= "001000";
					when "011000100110111" => rgb <= "001000";
					when "011000100111000" => rgb <= "001000";
					when "011000100111001" => rgb <= "001000";
					when "011000100111010" => rgb <= "001000";
					when "011000100111011" => rgb <= "001000";
					when "011000100111100" => rgb <= "001000";
					when "011000100111101" => rgb <= "001000";
					when "011000100111110" => rgb <= "001000";
					when "011000100111111" => rgb <= "001000";
					when "011000101000000" => rgb <= "001000";
					when "011000101000001" => rgb <= "001000";
					when "011000101000010" => rgb <= "001000";
					when "011000101000011" => rgb <= "001000";
					when "011000101000100" => rgb <= "001000";
					when "011000101000101" => rgb <= "001000";
					when "011000101000110" => rgb <= "001000";
					when "011000101000111" => rgb <= "001000";
					when "011000101001000" => rgb <= "001000";
					when "011000101001001" => rgb <= "001000";
					when "011000101001010" => rgb <= "001000";
					when "011000101001011" => rgb <= "001000";
					when "011000101001100" => rgb <= "001000";
					when "011000101001101" => rgb <= "001000";
					when "011000101001110" => rgb <= "001000";
					when "011000101001111" => rgb <= "001000";
					when "011000101010000" => rgb <= "001000";
					when "011000101010001" => rgb <= "001000";
					when "011000101010010" => rgb <= "001000";
					when "011000101010011" => rgb <= "001000";
					when "011000101010100" => rgb <= "000000";
					when "011000101010101" => rgb <= "000000";
					when "011000101010110" => rgb <= "101111";
					when "011000101010111" => rgb <= "101111";
					when "011000101011000" => rgb <= "101111";
					when "011000101011001" => rgb <= "101111";
					when "011000101011010" => rgb <= "101111";
					when "011000101011011" => rgb <= "101111";
					when "011000101011100" => rgb <= "101111";
					when "011000101011101" => rgb <= "101111";
					when "011000101011110" => rgb <= "101111";
					when "011000101011111" => rgb <= "101111";
					when "011000101100000" => rgb <= "101111";
					when "011000101100001" => rgb <= "101111";
					when "011000101100010" => rgb <= "101111";
					when "011000101100011" => rgb <= "101111";
					when "011000101100100" => rgb <= "101111";
					when "011000101100101" => rgb <= "101111";
					when "011000101100110" => rgb <= "101111";
					when "011000101100111" => rgb <= "101111";
					when "011000101101000" => rgb <= "101111";
					when "011000101101001" => rgb <= "101111";
					when "011000101101010" => rgb <= "101111";
					when "011000101101011" => rgb <= "101111";
					when "011000101101100" => rgb <= "101111";
					when "011000101101101" => rgb <= "101111";
					when "011000101101110" => rgb <= "101111";
					when "011000101101111" => rgb <= "101111";
					when "011000101110000" => rgb <= "101111";
					when "011000101110001" => rgb <= "101111";
					when "011000101110010" => rgb <= "101111";
					when "011000101110011" => rgb <= "101111";
					when "011000101110100" => rgb <= "101111";
					when "011000101110101" => rgb <= "101111";
					when "011000101110110" => rgb <= "101111";
					when "011000101110111" => rgb <= "101111";
					when "011000101111000" => rgb <= "101111";
					when "011000101111001" => rgb <= "101111";
					when "011000101111010" => rgb <= "101111";
					when "011000101111011" => rgb <= "101111";
					when "011000101111100" => rgb <= "101111";
					when "011000101111101" => rgb <= "101111";
					when "011000101111110" => rgb <= "101111";
					when "011000101111111" => rgb <= "101111";
					when "011000110000000" => rgb <= "101111";
					when "011000110000001" => rgb <= "101111";
					when "011000110000010" => rgb <= "101111";
					when "011000110000011" => rgb <= "101111";
					when "011000110000100" => rgb <= "101111";
					when "011000110000101" => rgb <= "101111";
					when "011000110000110" => rgb <= "101111";
					when "011000110000111" => rgb <= "101111";
					when "011000110001000" => rgb <= "101111";
					when "011000110001001" => rgb <= "101111";
					when "011000110001010" => rgb <= "101111";
					when "011000110001011" => rgb <= "101111";
					when "011000110001100" => rgb <= "101111";
					when "011000110001101" => rgb <= "101111";
					when "011000110001110" => rgb <= "101111";
					when "011000110001111" => rgb <= "101111";
					when "011000110010000" => rgb <= "101111";
					when "011000110010001" => rgb <= "101111";
					when "011000110010010" => rgb <= "101111";
					when "011000110010011" => rgb <= "101111";
					when "011000110010100" => rgb <= "101111";
					when "011000110010101" => rgb <= "101111";
					when "011000110010110" => rgb <= "101111";
					when "011000110010111" => rgb <= "101111";
					when "011000110011000" => rgb <= "101111";
					when "011000110011001" => rgb <= "101111";
					when "011000110011010" => rgb <= "101111";
					when "011000110011011" => rgb <= "101111";
					when "011000110011100" => rgb <= "101111";
					when "011000110011101" => rgb <= "101111";
					when "011000110011110" => rgb <= "101111";
					when "011000110011111" => rgb <= "101111";
					when "011001000000000" => rgb <= "001000";
					when "011001000000001" => rgb <= "001000";
					when "011001000000010" => rgb <= "001000";
					when "011001000000011" => rgb <= "001000";
					when "011001000000100" => rgb <= "001000";
					when "011001000000101" => rgb <= "001000";
					when "011001000000110" => rgb <= "001000";
					when "011001000000111" => rgb <= "001000";
					when "011001000001000" => rgb <= "001000";
					when "011001000001001" => rgb <= "001000";
					when "011001000001010" => rgb <= "001000";
					when "011001000001011" => rgb <= "001000";
					when "011001000001100" => rgb <= "001000";
					when "011001000001101" => rgb <= "001000";
					when "011001000001110" => rgb <= "001000";
					when "011001000001111" => rgb <= "001000";
					when "011001000010000" => rgb <= "001000";
					when "011001000010001" => rgb <= "001000";
					when "011001000010010" => rgb <= "001000";
					when "011001000010011" => rgb <= "001000";
					when "011001000010100" => rgb <= "001000";
					when "011001000010101" => rgb <= "001000";
					when "011001000010110" => rgb <= "001000";
					when "011001000010111" => rgb <= "001000";
					when "011001000011000" => rgb <= "001000";
					when "011001000011001" => rgb <= "001000";
					when "011001000011010" => rgb <= "001000";
					when "011001000011011" => rgb <= "001000";
					when "011001000011100" => rgb <= "001000";
					when "011001000011101" => rgb <= "001000";
					when "011001000011110" => rgb <= "001000";
					when "011001000011111" => rgb <= "001000";
					when "011001000100000" => rgb <= "001000";
					when "011001000100001" => rgb <= "001000";
					when "011001000100010" => rgb <= "001000";
					when "011001000100011" => rgb <= "001000";
					when "011001000100100" => rgb <= "001000";
					when "011001000100101" => rgb <= "001000";
					when "011001000100110" => rgb <= "001000";
					when "011001000100111" => rgb <= "001000";
					when "011001000101000" => rgb <= "001000";
					when "011001000101001" => rgb <= "001000";
					when "011001000101010" => rgb <= "001000";
					when "011001000101011" => rgb <= "001000";
					when "011001000101100" => rgb <= "001000";
					when "011001000101101" => rgb <= "001000";
					when "011001000101110" => rgb <= "001000";
					when "011001000101111" => rgb <= "001000";
					when "011001000110000" => rgb <= "001000";
					when "011001000110001" => rgb <= "001000";
					when "011001000110010" => rgb <= "001000";
					when "011001000110011" => rgb <= "001000";
					when "011001000110100" => rgb <= "001000";
					when "011001000110101" => rgb <= "001000";
					when "011001000110110" => rgb <= "001000";
					when "011001000110111" => rgb <= "001000";
					when "011001000111000" => rgb <= "001000";
					when "011001000111001" => rgb <= "001000";
					when "011001000111010" => rgb <= "001000";
					when "011001000111011" => rgb <= "001000";
					when "011001000111100" => rgb <= "001000";
					when "011001000111101" => rgb <= "001000";
					when "011001000111110" => rgb <= "001000";
					when "011001000111111" => rgb <= "001000";
					when "011001001000000" => rgb <= "001000";
					when "011001001000001" => rgb <= "001000";
					when "011001001000010" => rgb <= "001000";
					when "011001001000011" => rgb <= "001000";
					when "011001001000100" => rgb <= "001000";
					when "011001001000101" => rgb <= "001000";
					when "011001001000110" => rgb <= "001000";
					when "011001001000111" => rgb <= "001000";
					when "011001001001000" => rgb <= "001000";
					when "011001001001001" => rgb <= "001000";
					when "011001001001010" => rgb <= "001000";
					when "011001001001011" => rgb <= "001000";
					when "011001001001100" => rgb <= "001000";
					when "011001001001101" => rgb <= "001000";
					when "011001001001110" => rgb <= "001000";
					when "011001001001111" => rgb <= "001000";
					when "011001001010000" => rgb <= "001000";
					when "011001001010001" => rgb <= "001000";
					when "011001001010010" => rgb <= "001000";
					when "011001001010011" => rgb <= "001000";
					when "011001001010100" => rgb <= "001000";
					when "011001001010101" => rgb <= "001000";
					when "011001001010110" => rgb <= "000000";
					when "011001001010111" => rgb <= "000000";
					when "011001001011000" => rgb <= "101111";
					when "011001001011001" => rgb <= "101111";
					when "011001001011010" => rgb <= "101111";
					when "011001001011011" => rgb <= "101111";
					when "011001001011100" => rgb <= "101111";
					when "011001001011101" => rgb <= "101111";
					when "011001001011110" => rgb <= "101111";
					when "011001001011111" => rgb <= "101111";
					when "011001001100000" => rgb <= "101111";
					when "011001001100001" => rgb <= "101111";
					when "011001001100010" => rgb <= "101111";
					when "011001001100011" => rgb <= "101111";
					when "011001001100100" => rgb <= "101111";
					when "011001001100101" => rgb <= "101111";
					when "011001001100110" => rgb <= "101111";
					when "011001001100111" => rgb <= "101111";
					when "011001001101000" => rgb <= "101111";
					when "011001001101001" => rgb <= "101111";
					when "011001001101010" => rgb <= "101111";
					when "011001001101011" => rgb <= "101111";
					when "011001001101100" => rgb <= "101111";
					when "011001001101101" => rgb <= "101111";
					when "011001001101110" => rgb <= "101111";
					when "011001001101111" => rgb <= "101111";
					when "011001001110000" => rgb <= "101111";
					when "011001001110001" => rgb <= "101111";
					when "011001001110010" => rgb <= "101111";
					when "011001001110011" => rgb <= "101111";
					when "011001001110100" => rgb <= "101111";
					when "011001001110101" => rgb <= "101111";
					when "011001001110110" => rgb <= "101111";
					when "011001001110111" => rgb <= "101111";
					when "011001001111000" => rgb <= "101111";
					when "011001001111001" => rgb <= "101111";
					when "011001001111010" => rgb <= "101111";
					when "011001001111011" => rgb <= "101111";
					when "011001001111100" => rgb <= "101111";
					when "011001001111101" => rgb <= "101111";
					when "011001001111110" => rgb <= "101111";
					when "011001001111111" => rgb <= "101111";
					when "011001010000000" => rgb <= "101111";
					when "011001010000001" => rgb <= "101111";
					when "011001010000010" => rgb <= "101111";
					when "011001010000011" => rgb <= "101111";
					when "011001010000100" => rgb <= "101111";
					when "011001010000101" => rgb <= "101111";
					when "011001010000110" => rgb <= "101111";
					when "011001010000111" => rgb <= "101111";
					when "011001010001000" => rgb <= "101111";
					when "011001010001001" => rgb <= "101111";
					when "011001010001010" => rgb <= "101111";
					when "011001010001011" => rgb <= "101111";
					when "011001010001100" => rgb <= "101111";
					when "011001010001101" => rgb <= "101111";
					when "011001010001110" => rgb <= "101111";
					when "011001010001111" => rgb <= "101111";
					when "011001010010000" => rgb <= "101111";
					when "011001010010001" => rgb <= "101111";
					when "011001010010010" => rgb <= "101111";
					when "011001010010011" => rgb <= "101111";
					when "011001010010100" => rgb <= "101111";
					when "011001010010101" => rgb <= "101111";
					when "011001010010110" => rgb <= "101111";
					when "011001010010111" => rgb <= "101111";
					when "011001010011000" => rgb <= "101111";
					when "011001010011001" => rgb <= "101111";
					when "011001010011010" => rgb <= "101111";
					when "011001010011011" => rgb <= "101111";
					when "011001010011100" => rgb <= "101111";
					when "011001010011101" => rgb <= "101111";
					when "011001010011110" => rgb <= "101111";
					when "011001010011111" => rgb <= "101111";
					when "011001100000000" => rgb <= "001000";
					when "011001100000001" => rgb <= "001000";
					when "011001100000010" => rgb <= "001000";
					when "011001100000011" => rgb <= "001000";
					when "011001100000100" => rgb <= "001000";
					when "011001100000101" => rgb <= "001000";
					when "011001100000110" => rgb <= "001000";
					when "011001100000111" => rgb <= "001000";
					when "011001100001000" => rgb <= "001000";
					when "011001100001001" => rgb <= "001000";
					when "011001100001010" => rgb <= "001000";
					when "011001100001011" => rgb <= "001000";
					when "011001100001100" => rgb <= "001000";
					when "011001100001101" => rgb <= "001000";
					when "011001100001110" => rgb <= "001000";
					when "011001100001111" => rgb <= "001000";
					when "011001100010000" => rgb <= "001000";
					when "011001100010001" => rgb <= "001000";
					when "011001100010010" => rgb <= "001000";
					when "011001100010011" => rgb <= "001000";
					when "011001100010100" => rgb <= "001000";
					when "011001100010101" => rgb <= "001000";
					when "011001100010110" => rgb <= "001000";
					when "011001100010111" => rgb <= "001000";
					when "011001100011000" => rgb <= "001000";
					when "011001100011001" => rgb <= "001000";
					when "011001100011010" => rgb <= "001000";
					when "011001100011011" => rgb <= "001000";
					when "011001100011100" => rgb <= "001000";
					when "011001100011101" => rgb <= "001000";
					when "011001100011110" => rgb <= "001000";
					when "011001100011111" => rgb <= "001000";
					when "011001100100000" => rgb <= "001000";
					when "011001100100001" => rgb <= "001000";
					when "011001100100010" => rgb <= "001000";
					when "011001100100011" => rgb <= "001000";
					when "011001100100100" => rgb <= "001000";
					when "011001100100101" => rgb <= "001000";
					when "011001100100110" => rgb <= "001000";
					when "011001100100111" => rgb <= "001000";
					when "011001100101000" => rgb <= "001000";
					when "011001100101001" => rgb <= "001000";
					when "011001100101010" => rgb <= "001000";
					when "011001100101011" => rgb <= "001000";
					when "011001100101100" => rgb <= "001000";
					when "011001100101101" => rgb <= "001000";
					when "011001100101110" => rgb <= "001000";
					when "011001100101111" => rgb <= "001000";
					when "011001100110000" => rgb <= "001000";
					when "011001100110001" => rgb <= "001000";
					when "011001100110010" => rgb <= "001000";
					when "011001100110011" => rgb <= "001000";
					when "011001100110100" => rgb <= "001000";
					when "011001100110101" => rgb <= "001000";
					when "011001100110110" => rgb <= "001000";
					when "011001100110111" => rgb <= "001000";
					when "011001100111000" => rgb <= "001000";
					when "011001100111001" => rgb <= "001000";
					when "011001100111010" => rgb <= "001000";
					when "011001100111011" => rgb <= "001000";
					when "011001100111100" => rgb <= "001000";
					when "011001100111101" => rgb <= "001000";
					when "011001100111110" => rgb <= "001000";
					when "011001100111111" => rgb <= "001000";
					when "011001101000000" => rgb <= "001000";
					when "011001101000001" => rgb <= "001000";
					when "011001101000010" => rgb <= "001000";
					when "011001101000011" => rgb <= "001000";
					when "011001101000100" => rgb <= "001000";
					when "011001101000101" => rgb <= "001000";
					when "011001101000110" => rgb <= "001000";
					when "011001101000111" => rgb <= "001000";
					when "011001101001000" => rgb <= "001000";
					when "011001101001001" => rgb <= "001000";
					when "011001101001010" => rgb <= "001000";
					when "011001101001011" => rgb <= "001000";
					when "011001101001100" => rgb <= "001000";
					when "011001101001101" => rgb <= "001000";
					when "011001101001110" => rgb <= "001000";
					when "011001101001111" => rgb <= "001000";
					when "011001101010000" => rgb <= "001000";
					when "011001101010001" => rgb <= "001000";
					when "011001101010010" => rgb <= "001000";
					when "011001101010011" => rgb <= "001000";
					when "011001101010100" => rgb <= "001000";
					when "011001101010101" => rgb <= "001000";
					when "011001101010110" => rgb <= "000000";
					when "011001101010111" => rgb <= "000000";
					when "011001101011000" => rgb <= "101111";
					when "011001101011001" => rgb <= "101111";
					when "011001101011010" => rgb <= "101111";
					when "011001101011011" => rgb <= "101111";
					when "011001101011100" => rgb <= "101111";
					when "011001101011101" => rgb <= "101111";
					when "011001101011110" => rgb <= "101111";
					when "011001101011111" => rgb <= "101111";
					when "011001101100000" => rgb <= "101111";
					when "011001101100001" => rgb <= "101111";
					when "011001101100010" => rgb <= "101111";
					when "011001101100011" => rgb <= "101111";
					when "011001101100100" => rgb <= "101111";
					when "011001101100101" => rgb <= "101111";
					when "011001101100110" => rgb <= "101111";
					when "011001101100111" => rgb <= "101111";
					when "011001101101000" => rgb <= "101111";
					when "011001101101001" => rgb <= "101111";
					when "011001101101010" => rgb <= "101111";
					when "011001101101011" => rgb <= "101111";
					when "011001101101100" => rgb <= "101111";
					when "011001101101101" => rgb <= "101111";
					when "011001101101110" => rgb <= "101111";
					when "011001101101111" => rgb <= "101111";
					when "011001101110000" => rgb <= "101111";
					when "011001101110001" => rgb <= "101111";
					when "011001101110010" => rgb <= "101111";
					when "011001101110011" => rgb <= "101111";
					when "011001101110100" => rgb <= "101111";
					when "011001101110101" => rgb <= "101111";
					when "011001101110110" => rgb <= "101111";
					when "011001101110111" => rgb <= "101111";
					when "011001101111000" => rgb <= "101111";
					when "011001101111001" => rgb <= "101111";
					when "011001101111010" => rgb <= "101111";
					when "011001101111011" => rgb <= "101111";
					when "011001101111100" => rgb <= "101111";
					when "011001101111101" => rgb <= "101111";
					when "011001101111110" => rgb <= "101111";
					when "011001101111111" => rgb <= "101111";
					when "011001110000000" => rgb <= "101111";
					when "011001110000001" => rgb <= "101111";
					when "011001110000010" => rgb <= "101111";
					when "011001110000011" => rgb <= "101111";
					when "011001110000100" => rgb <= "101111";
					when "011001110000101" => rgb <= "101111";
					when "011001110000110" => rgb <= "101111";
					when "011001110000111" => rgb <= "101111";
					when "011001110001000" => rgb <= "101111";
					when "011001110001001" => rgb <= "101111";
					when "011001110001010" => rgb <= "101111";
					when "011001110001011" => rgb <= "101111";
					when "011001110001100" => rgb <= "101111";
					when "011001110001101" => rgb <= "101111";
					when "011001110001110" => rgb <= "101111";
					when "011001110001111" => rgb <= "101111";
					when "011001110010000" => rgb <= "101111";
					when "011001110010001" => rgb <= "101111";
					when "011001110010010" => rgb <= "101111";
					when "011001110010011" => rgb <= "101111";
					when "011001110010100" => rgb <= "101111";
					when "011001110010101" => rgb <= "101111";
					when "011001110010110" => rgb <= "101111";
					when "011001110010111" => rgb <= "101111";
					when "011001110011000" => rgb <= "101111";
					when "011001110011001" => rgb <= "101111";
					when "011001110011010" => rgb <= "101111";
					when "011001110011011" => rgb <= "101111";
					when "011001110011100" => rgb <= "101111";
					when "011001110011101" => rgb <= "101111";
					when "011001110011110" => rgb <= "101111";
					when "011001110011111" => rgb <= "101111";
					when "011010000000000" => rgb <= "001000";
					when "011010000000001" => rgb <= "001000";
					when "011010000000010" => rgb <= "001000";
					when "011010000000011" => rgb <= "001000";
					when "011010000000100" => rgb <= "001000";
					when "011010000000101" => rgb <= "001000";
					when "011010000000110" => rgb <= "001000";
					when "011010000000111" => rgb <= "001000";
					when "011010000001000" => rgb <= "001000";
					when "011010000001001" => rgb <= "001000";
					when "011010000001010" => rgb <= "001000";
					when "011010000001011" => rgb <= "001000";
					when "011010000001100" => rgb <= "001000";
					when "011010000001101" => rgb <= "001000";
					when "011010000001110" => rgb <= "001000";
					when "011010000001111" => rgb <= "001000";
					when "011010000010000" => rgb <= "001000";
					when "011010000010001" => rgb <= "001000";
					when "011010000010010" => rgb <= "001000";
					when "011010000010011" => rgb <= "001000";
					when "011010000010100" => rgb <= "001000";
					when "011010000010101" => rgb <= "001000";
					when "011010000010110" => rgb <= "001000";
					when "011010000010111" => rgb <= "001000";
					when "011010000011000" => rgb <= "001000";
					when "011010000011001" => rgb <= "001000";
					when "011010000011010" => rgb <= "001000";
					when "011010000011011" => rgb <= "001000";
					when "011010000011100" => rgb <= "001000";
					when "011010000011101" => rgb <= "001000";
					when "011010000011110" => rgb <= "001000";
					when "011010000011111" => rgb <= "001000";
					when "011010000100000" => rgb <= "001000";
					when "011010000100001" => rgb <= "001000";
					when "011010000100010" => rgb <= "001000";
					when "011010000100011" => rgb <= "001000";
					when "011010000100100" => rgb <= "001000";
					when "011010000100101" => rgb <= "001000";
					when "011010000100110" => rgb <= "001000";
					when "011010000100111" => rgb <= "001000";
					when "011010000101000" => rgb <= "001000";
					when "011010000101001" => rgb <= "001000";
					when "011010000101010" => rgb <= "001000";
					when "011010000101011" => rgb <= "001000";
					when "011010000101100" => rgb <= "001000";
					when "011010000101101" => rgb <= "001000";
					when "011010000101110" => rgb <= "001000";
					when "011010000101111" => rgb <= "001000";
					when "011010000110000" => rgb <= "001000";
					when "011010000110001" => rgb <= "001000";
					when "011010000110010" => rgb <= "001000";
					when "011010000110011" => rgb <= "001000";
					when "011010000110100" => rgb <= "001000";
					when "011010000110101" => rgb <= "001000";
					when "011010000110110" => rgb <= "001000";
					when "011010000110111" => rgb <= "001000";
					when "011010000111000" => rgb <= "001000";
					when "011010000111001" => rgb <= "001000";
					when "011010000111010" => rgb <= "001000";
					when "011010000111011" => rgb <= "001000";
					when "011010000111100" => rgb <= "001000";
					when "011010000111101" => rgb <= "001000";
					when "011010000111110" => rgb <= "001000";
					when "011010000111111" => rgb <= "001000";
					when "011010001000000" => rgb <= "001000";
					when "011010001000001" => rgb <= "001000";
					when "011010001000010" => rgb <= "001000";
					when "011010001000011" => rgb <= "001000";
					when "011010001000100" => rgb <= "001000";
					when "011010001000101" => rgb <= "001000";
					when "011010001000110" => rgb <= "001000";
					when "011010001000111" => rgb <= "001000";
					when "011010001001000" => rgb <= "001000";
					when "011010001001001" => rgb <= "001000";
					when "011010001001010" => rgb <= "001000";
					when "011010001001011" => rgb <= "001000";
					when "011010001001100" => rgb <= "001000";
					when "011010001001101" => rgb <= "001000";
					when "011010001001110" => rgb <= "001000";
					when "011010001001111" => rgb <= "001000";
					when "011010001010000" => rgb <= "001000";
					when "011010001010001" => rgb <= "001000";
					when "011010001010010" => rgb <= "001000";
					when "011010001010011" => rgb <= "001000";
					when "011010001010100" => rgb <= "001000";
					when "011010001010101" => rgb <= "001000";
					when "011010001010110" => rgb <= "000000";
					when "011010001010111" => rgb <= "000000";
					when "011010001011000" => rgb <= "101111";
					when "011010001011001" => rgb <= "101111";
					when "011010001011010" => rgb <= "101111";
					when "011010001011011" => rgb <= "101111";
					when "011010001011100" => rgb <= "101111";
					when "011010001011101" => rgb <= "101111";
					when "011010001011110" => rgb <= "101111";
					when "011010001011111" => rgb <= "101111";
					when "011010001100000" => rgb <= "101111";
					when "011010001100001" => rgb <= "101111";
					when "011010001100010" => rgb <= "101111";
					when "011010001100011" => rgb <= "101111";
					when "011010001100100" => rgb <= "101111";
					when "011010001100101" => rgb <= "101111";
					when "011010001100110" => rgb <= "101111";
					when "011010001100111" => rgb <= "101111";
					when "011010001101000" => rgb <= "101111";
					when "011010001101001" => rgb <= "101111";
					when "011010001101010" => rgb <= "101111";
					when "011010001101011" => rgb <= "101111";
					when "011010001101100" => rgb <= "101111";
					when "011010001101101" => rgb <= "101111";
					when "011010001101110" => rgb <= "101111";
					when "011010001101111" => rgb <= "101111";
					when "011010001110000" => rgb <= "101111";
					when "011010001110001" => rgb <= "101111";
					when "011010001110010" => rgb <= "101111";
					when "011010001110011" => rgb <= "101111";
					when "011010001110100" => rgb <= "101111";
					when "011010001110101" => rgb <= "101111";
					when "011010001110110" => rgb <= "101111";
					when "011010001110111" => rgb <= "101111";
					when "011010001111000" => rgb <= "101111";
					when "011010001111001" => rgb <= "101111";
					when "011010001111010" => rgb <= "101111";
					when "011010001111011" => rgb <= "101111";
					when "011010001111100" => rgb <= "101111";
					when "011010001111101" => rgb <= "101111";
					when "011010001111110" => rgb <= "101111";
					when "011010001111111" => rgb <= "101111";
					when "011010010000000" => rgb <= "101111";
					when "011010010000001" => rgb <= "101111";
					when "011010010000010" => rgb <= "101111";
					when "011010010000011" => rgb <= "101111";
					when "011010010000100" => rgb <= "101111";
					when "011010010000101" => rgb <= "101111";
					when "011010010000110" => rgb <= "101111";
					when "011010010000111" => rgb <= "101111";
					when "011010010001000" => rgb <= "101111";
					when "011010010001001" => rgb <= "101111";
					when "011010010001010" => rgb <= "101111";
					when "011010010001011" => rgb <= "101111";
					when "011010010001100" => rgb <= "101111";
					when "011010010001101" => rgb <= "101111";
					when "011010010001110" => rgb <= "101111";
					when "011010010001111" => rgb <= "101111";
					when "011010010010000" => rgb <= "101111";
					when "011010010010001" => rgb <= "101111";
					when "011010010010010" => rgb <= "101111";
					when "011010010010011" => rgb <= "101111";
					when "011010010010100" => rgb <= "101111";
					when "011010010010101" => rgb <= "101111";
					when "011010010010110" => rgb <= "101111";
					when "011010010010111" => rgb <= "101111";
					when "011010010011000" => rgb <= "101111";
					when "011010010011001" => rgb <= "101111";
					when "011010010011010" => rgb <= "101111";
					when "011010010011011" => rgb <= "101111";
					when "011010010011100" => rgb <= "101111";
					when "011010010011101" => rgb <= "101111";
					when "011010010011110" => rgb <= "101111";
					when "011010010011111" => rgb <= "101111";
					when "011010100000000" => rgb <= "001000";
					when "011010100000001" => rgb <= "001000";
					when "011010100000010" => rgb <= "001000";
					when "011010100000011" => rgb <= "001000";
					when "011010100000100" => rgb <= "001000";
					when "011010100000101" => rgb <= "001000";
					when "011010100000110" => rgb <= "001000";
					when "011010100000111" => rgb <= "001000";
					when "011010100001000" => rgb <= "001000";
					when "011010100001001" => rgb <= "001000";
					when "011010100001010" => rgb <= "001000";
					when "011010100001011" => rgb <= "001000";
					when "011010100001100" => rgb <= "001000";
					when "011010100001101" => rgb <= "001000";
					when "011010100001110" => rgb <= "001000";
					when "011010100001111" => rgb <= "001000";
					when "011010100010000" => rgb <= "001000";
					when "011010100010001" => rgb <= "001000";
					when "011010100010010" => rgb <= "001000";
					when "011010100010011" => rgb <= "001000";
					when "011010100010100" => rgb <= "001000";
					when "011010100010101" => rgb <= "001000";
					when "011010100010110" => rgb <= "001000";
					when "011010100010111" => rgb <= "001000";
					when "011010100011000" => rgb <= "001000";
					when "011010100011001" => rgb <= "001000";
					when "011010100011010" => rgb <= "001000";
					when "011010100011011" => rgb <= "001000";
					when "011010100011100" => rgb <= "001000";
					when "011010100011101" => rgb <= "001000";
					when "011010100011110" => rgb <= "001000";
					when "011010100011111" => rgb <= "001000";
					when "011010100100000" => rgb <= "001000";
					when "011010100100001" => rgb <= "001000";
					when "011010100100010" => rgb <= "001000";
					when "011010100100011" => rgb <= "001000";
					when "011010100100100" => rgb <= "001000";
					when "011010100100101" => rgb <= "001000";
					when "011010100100110" => rgb <= "001000";
					when "011010100100111" => rgb <= "001000";
					when "011010100101000" => rgb <= "001000";
					when "011010100101001" => rgb <= "001000";
					when "011010100101010" => rgb <= "001000";
					when "011010100101011" => rgb <= "001000";
					when "011010100101100" => rgb <= "001000";
					when "011010100101101" => rgb <= "001000";
					when "011010100101110" => rgb <= "001000";
					when "011010100101111" => rgb <= "001000";
					when "011010100110000" => rgb <= "001000";
					when "011010100110001" => rgb <= "001000";
					when "011010100110010" => rgb <= "001000";
					when "011010100110011" => rgb <= "001000";
					when "011010100110100" => rgb <= "001000";
					when "011010100110101" => rgb <= "001000";
					when "011010100110110" => rgb <= "001000";
					when "011010100110111" => rgb <= "001000";
					when "011010100111000" => rgb <= "001000";
					when "011010100111001" => rgb <= "001000";
					when "011010100111010" => rgb <= "001000";
					when "011010100111011" => rgb <= "001000";
					when "011010100111100" => rgb <= "001000";
					when "011010100111101" => rgb <= "001000";
					when "011010100111110" => rgb <= "001000";
					when "011010100111111" => rgb <= "001000";
					when "011010101000000" => rgb <= "001000";
					when "011010101000001" => rgb <= "001000";
					when "011010101000010" => rgb <= "001000";
					when "011010101000011" => rgb <= "001000";
					when "011010101000100" => rgb <= "001000";
					when "011010101000101" => rgb <= "001000";
					when "011010101000110" => rgb <= "001000";
					when "011010101000111" => rgb <= "001000";
					when "011010101001000" => rgb <= "001000";
					when "011010101001001" => rgb <= "001000";
					when "011010101001010" => rgb <= "001000";
					when "011010101001011" => rgb <= "001000";
					when "011010101001100" => rgb <= "001000";
					when "011010101001101" => rgb <= "001000";
					when "011010101001110" => rgb <= "001000";
					when "011010101001111" => rgb <= "001000";
					when "011010101010000" => rgb <= "001000";
					when "011010101010001" => rgb <= "001000";
					when "011010101010010" => rgb <= "001000";
					when "011010101010011" => rgb <= "001000";
					when "011010101010100" => rgb <= "001000";
					when "011010101010101" => rgb <= "001000";
					when "011010101010110" => rgb <= "000000";
					when "011010101010111" => rgb <= "000000";
					when "011010101011000" => rgb <= "101111";
					when "011010101011001" => rgb <= "101111";
					when "011010101011010" => rgb <= "101111";
					when "011010101011011" => rgb <= "101111";
					when "011010101011100" => rgb <= "101111";
					when "011010101011101" => rgb <= "101111";
					when "011010101011110" => rgb <= "101111";
					when "011010101011111" => rgb <= "101111";
					when "011010101100000" => rgb <= "101111";
					when "011010101100001" => rgb <= "101111";
					when "011010101100010" => rgb <= "101111";
					when "011010101100011" => rgb <= "101111";
					when "011010101100100" => rgb <= "101111";
					when "011010101100101" => rgb <= "101111";
					when "011010101100110" => rgb <= "101111";
					when "011010101100111" => rgb <= "101111";
					when "011010101101000" => rgb <= "101111";
					when "011010101101001" => rgb <= "101111";
					when "011010101101010" => rgb <= "101111";
					when "011010101101011" => rgb <= "101111";
					when "011010101101100" => rgb <= "101111";
					when "011010101101101" => rgb <= "101111";
					when "011010101101110" => rgb <= "101111";
					when "011010101101111" => rgb <= "101111";
					when "011010101110000" => rgb <= "101111";
					when "011010101110001" => rgb <= "101111";
					when "011010101110010" => rgb <= "101111";
					when "011010101110011" => rgb <= "101111";
					when "011010101110100" => rgb <= "101111";
					when "011010101110101" => rgb <= "101111";
					when "011010101110110" => rgb <= "101111";
					when "011010101110111" => rgb <= "101111";
					when "011010101111000" => rgb <= "101111";
					when "011010101111001" => rgb <= "101111";
					when "011010101111010" => rgb <= "101111";
					when "011010101111011" => rgb <= "101111";
					when "011010101111100" => rgb <= "101111";
					when "011010101111101" => rgb <= "101111";
					when "011010101111110" => rgb <= "101111";
					when "011010101111111" => rgb <= "101111";
					when "011010110000000" => rgb <= "101111";
					when "011010110000001" => rgb <= "101111";
					when "011010110000010" => rgb <= "101111";
					when "011010110000011" => rgb <= "101111";
					when "011010110000100" => rgb <= "101111";
					when "011010110000101" => rgb <= "101111";
					when "011010110000110" => rgb <= "101111";
					when "011010110000111" => rgb <= "101111";
					when "011010110001000" => rgb <= "101111";
					when "011010110001001" => rgb <= "101111";
					when "011010110001010" => rgb <= "101111";
					when "011010110001011" => rgb <= "101111";
					when "011010110001100" => rgb <= "101111";
					when "011010110001101" => rgb <= "101111";
					when "011010110001110" => rgb <= "101111";
					when "011010110001111" => rgb <= "101111";
					when "011010110010000" => rgb <= "101111";
					when "011010110010001" => rgb <= "101111";
					when "011010110010010" => rgb <= "101111";
					when "011010110010011" => rgb <= "101111";
					when "011010110010100" => rgb <= "101111";
					when "011010110010101" => rgb <= "101111";
					when "011010110010110" => rgb <= "101111";
					when "011010110010111" => rgb <= "101111";
					when "011010110011000" => rgb <= "101111";
					when "011010110011001" => rgb <= "101111";
					when "011010110011010" => rgb <= "101111";
					when "011010110011011" => rgb <= "101111";
					when "011010110011100" => rgb <= "101111";
					when "011010110011101" => rgb <= "101111";
					when "011010110011110" => rgb <= "101111";
					when "011010110011111" => rgb <= "101111";
					when "011011000000000" => rgb <= "001000";
					when "011011000000001" => rgb <= "001000";
					when "011011000000010" => rgb <= "001000";
					when "011011000000011" => rgb <= "001000";
					when "011011000000100" => rgb <= "001000";
					when "011011000000101" => rgb <= "001000";
					when "011011000000110" => rgb <= "001000";
					when "011011000000111" => rgb <= "001000";
					when "011011000001000" => rgb <= "001000";
					when "011011000001001" => rgb <= "001000";
					when "011011000001010" => rgb <= "001000";
					when "011011000001011" => rgb <= "001000";
					when "011011000001100" => rgb <= "001000";
					when "011011000001101" => rgb <= "001000";
					when "011011000001110" => rgb <= "001000";
					when "011011000001111" => rgb <= "001000";
					when "011011000010000" => rgb <= "001000";
					when "011011000010001" => rgb <= "001000";
					when "011011000010010" => rgb <= "001000";
					when "011011000010011" => rgb <= "001000";
					when "011011000010100" => rgb <= "001000";
					when "011011000010101" => rgb <= "001000";
					when "011011000010110" => rgb <= "001000";
					when "011011000010111" => rgb <= "001000";
					when "011011000011000" => rgb <= "001000";
					when "011011000011001" => rgb <= "001000";
					when "011011000011010" => rgb <= "001000";
					when "011011000011011" => rgb <= "001000";
					when "011011000011100" => rgb <= "001000";
					when "011011000011101" => rgb <= "001000";
					when "011011000011110" => rgb <= "001000";
					when "011011000011111" => rgb <= "001000";
					when "011011000100000" => rgb <= "001000";
					when "011011000100001" => rgb <= "001000";
					when "011011000100010" => rgb <= "001000";
					when "011011000100011" => rgb <= "001000";
					when "011011000100100" => rgb <= "001000";
					when "011011000100101" => rgb <= "001000";
					when "011011000100110" => rgb <= "001000";
					when "011011000100111" => rgb <= "001000";
					when "011011000101000" => rgb <= "001000";
					when "011011000101001" => rgb <= "001000";
					when "011011000101010" => rgb <= "001000";
					when "011011000101011" => rgb <= "001000";
					when "011011000101100" => rgb <= "001000";
					when "011011000101101" => rgb <= "001000";
					when "011011000101110" => rgb <= "001000";
					when "011011000101111" => rgb <= "001000";
					when "011011000110000" => rgb <= "001000";
					when "011011000110001" => rgb <= "001000";
					when "011011000110010" => rgb <= "001000";
					when "011011000110011" => rgb <= "001000";
					when "011011000110100" => rgb <= "001000";
					when "011011000110101" => rgb <= "001000";
					when "011011000110110" => rgb <= "001000";
					when "011011000110111" => rgb <= "001000";
					when "011011000111000" => rgb <= "001000";
					when "011011000111001" => rgb <= "001000";
					when "011011000111010" => rgb <= "001000";
					when "011011000111011" => rgb <= "001000";
					when "011011000111100" => rgb <= "001000";
					when "011011000111101" => rgb <= "001000";
					when "011011000111110" => rgb <= "001000";
					when "011011000111111" => rgb <= "001000";
					when "011011001000000" => rgb <= "001000";
					when "011011001000001" => rgb <= "001000";
					when "011011001000010" => rgb <= "001000";
					when "011011001000011" => rgb <= "001000";
					when "011011001000100" => rgb <= "001000";
					when "011011001000101" => rgb <= "001000";
					when "011011001000110" => rgb <= "001000";
					when "011011001000111" => rgb <= "001000";
					when "011011001001000" => rgb <= "001000";
					when "011011001001001" => rgb <= "001000";
					when "011011001001010" => rgb <= "001000";
					when "011011001001011" => rgb <= "001000";
					when "011011001001100" => rgb <= "001000";
					when "011011001001101" => rgb <= "001000";
					when "011011001001110" => rgb <= "001000";
					when "011011001001111" => rgb <= "001000";
					when "011011001010000" => rgb <= "001000";
					when "011011001010001" => rgb <= "001000";
					when "011011001010010" => rgb <= "001000";
					when "011011001010011" => rgb <= "001000";
					when "011011001010100" => rgb <= "001000";
					when "011011001010101" => rgb <= "001000";
					when "011011001010110" => rgb <= "000000";
					when "011011001010111" => rgb <= "000000";
					when "011011001011000" => rgb <= "101111";
					when "011011001011001" => rgb <= "101111";
					when "011011001011010" => rgb <= "101111";
					when "011011001011011" => rgb <= "101111";
					when "011011001011100" => rgb <= "101111";
					when "011011001011101" => rgb <= "101111";
					when "011011001011110" => rgb <= "101111";
					when "011011001011111" => rgb <= "101111";
					when "011011001100000" => rgb <= "101111";
					when "011011001100001" => rgb <= "101111";
					when "011011001100010" => rgb <= "101111";
					when "011011001100011" => rgb <= "101111";
					when "011011001100100" => rgb <= "101111";
					when "011011001100101" => rgb <= "101111";
					when "011011001100110" => rgb <= "101111";
					when "011011001100111" => rgb <= "101111";
					when "011011001101000" => rgb <= "101111";
					when "011011001101001" => rgb <= "101111";
					when "011011001101010" => rgb <= "101111";
					when "011011001101011" => rgb <= "101111";
					when "011011001101100" => rgb <= "101111";
					when "011011001101101" => rgb <= "101111";
					when "011011001101110" => rgb <= "101111";
					when "011011001101111" => rgb <= "101111";
					when "011011001110000" => rgb <= "101111";
					when "011011001110001" => rgb <= "101111";
					when "011011001110010" => rgb <= "101111";
					when "011011001110011" => rgb <= "101111";
					when "011011001110100" => rgb <= "101111";
					when "011011001110101" => rgb <= "101111";
					when "011011001110110" => rgb <= "101111";
					when "011011001110111" => rgb <= "101111";
					when "011011001111000" => rgb <= "101111";
					when "011011001111001" => rgb <= "101111";
					when "011011001111010" => rgb <= "101111";
					when "011011001111011" => rgb <= "101111";
					when "011011001111100" => rgb <= "101111";
					when "011011001111101" => rgb <= "101111";
					when "011011001111110" => rgb <= "101111";
					when "011011001111111" => rgb <= "101111";
					when "011011010000000" => rgb <= "101111";
					when "011011010000001" => rgb <= "101111";
					when "011011010000010" => rgb <= "101111";
					when "011011010000011" => rgb <= "101111";
					when "011011010000100" => rgb <= "101111";
					when "011011010000101" => rgb <= "101111";
					when "011011010000110" => rgb <= "101111";
					when "011011010000111" => rgb <= "101111";
					when "011011010001000" => rgb <= "101111";
					when "011011010001001" => rgb <= "101111";
					when "011011010001010" => rgb <= "101111";
					when "011011010001011" => rgb <= "101111";
					when "011011010001100" => rgb <= "101111";
					when "011011010001101" => rgb <= "101111";
					when "011011010001110" => rgb <= "101111";
					when "011011010001111" => rgb <= "101111";
					when "011011010010000" => rgb <= "101111";
					when "011011010010001" => rgb <= "101111";
					when "011011010010010" => rgb <= "101111";
					when "011011010010011" => rgb <= "101111";
					when "011011010010100" => rgb <= "101111";
					when "011011010010101" => rgb <= "101111";
					when "011011010010110" => rgb <= "101111";
					when "011011010010111" => rgb <= "101111";
					when "011011010011000" => rgb <= "101111";
					when "011011010011001" => rgb <= "101111";
					when "011011010011010" => rgb <= "101111";
					when "011011010011011" => rgb <= "101111";
					when "011011010011100" => rgb <= "101111";
					when "011011010011101" => rgb <= "101111";
					when "011011010011110" => rgb <= "101111";
					when "011011010011111" => rgb <= "101111";
					when "011011100000000" => rgb <= "001000";
					when "011011100000001" => rgb <= "001000";
					when "011011100000010" => rgb <= "001000";
					when "011011100000011" => rgb <= "001000";
					when "011011100000100" => rgb <= "001000";
					when "011011100000101" => rgb <= "001000";
					when "011011100000110" => rgb <= "001000";
					when "011011100000111" => rgb <= "001000";
					when "011011100001000" => rgb <= "001000";
					when "011011100001001" => rgb <= "001000";
					when "011011100001010" => rgb <= "001000";
					when "011011100001011" => rgb <= "001000";
					when "011011100001100" => rgb <= "001000";
					when "011011100001101" => rgb <= "001000";
					when "011011100001110" => rgb <= "001000";
					when "011011100001111" => rgb <= "001000";
					when "011011100010000" => rgb <= "001000";
					when "011011100010001" => rgb <= "001000";
					when "011011100010010" => rgb <= "001000";
					when "011011100010011" => rgb <= "001000";
					when "011011100010100" => rgb <= "001000";
					when "011011100010101" => rgb <= "001000";
					when "011011100010110" => rgb <= "001000";
					when "011011100010111" => rgb <= "001000";
					when "011011100011000" => rgb <= "001000";
					when "011011100011001" => rgb <= "001000";
					when "011011100011010" => rgb <= "001000";
					when "011011100011011" => rgb <= "001000";
					when "011011100011100" => rgb <= "001000";
					when "011011100011101" => rgb <= "001000";
					when "011011100011110" => rgb <= "001000";
					when "011011100011111" => rgb <= "001000";
					when "011011100100000" => rgb <= "001000";
					when "011011100100001" => rgb <= "001000";
					when "011011100100010" => rgb <= "001000";
					when "011011100100011" => rgb <= "001000";
					when "011011100100100" => rgb <= "001000";
					when "011011100100101" => rgb <= "001000";
					when "011011100100110" => rgb <= "001000";
					when "011011100100111" => rgb <= "001000";
					when "011011100101000" => rgb <= "001000";
					when "011011100101001" => rgb <= "001000";
					when "011011100101010" => rgb <= "001000";
					when "011011100101011" => rgb <= "001000";
					when "011011100101100" => rgb <= "001000";
					when "011011100101101" => rgb <= "001000";
					when "011011100101110" => rgb <= "001000";
					when "011011100101111" => rgb <= "001000";
					when "011011100110000" => rgb <= "001000";
					when "011011100110001" => rgb <= "001000";
					when "011011100110010" => rgb <= "001000";
					when "011011100110011" => rgb <= "001000";
					when "011011100110100" => rgb <= "001000";
					when "011011100110101" => rgb <= "001000";
					when "011011100110110" => rgb <= "001000";
					when "011011100110111" => rgb <= "001000";
					when "011011100111000" => rgb <= "001000";
					when "011011100111001" => rgb <= "001000";
					when "011011100111010" => rgb <= "001000";
					when "011011100111011" => rgb <= "001000";
					when "011011100111100" => rgb <= "001000";
					when "011011100111101" => rgb <= "001000";
					when "011011100111110" => rgb <= "001000";
					when "011011100111111" => rgb <= "001000";
					when "011011101000000" => rgb <= "001000";
					when "011011101000001" => rgb <= "001000";
					when "011011101000010" => rgb <= "001000";
					when "011011101000011" => rgb <= "001000";
					when "011011101000100" => rgb <= "001000";
					when "011011101000101" => rgb <= "001000";
					when "011011101000110" => rgb <= "001000";
					when "011011101000111" => rgb <= "001000";
					when "011011101001000" => rgb <= "001000";
					when "011011101001001" => rgb <= "001000";
					when "011011101001010" => rgb <= "001000";
					when "011011101001011" => rgb <= "001000";
					when "011011101001100" => rgb <= "001000";
					when "011011101001101" => rgb <= "001000";
					when "011011101001110" => rgb <= "001000";
					when "011011101001111" => rgb <= "001000";
					when "011011101010000" => rgb <= "001000";
					when "011011101010001" => rgb <= "001000";
					when "011011101010010" => rgb <= "001000";
					when "011011101010011" => rgb <= "001000";
					when "011011101010100" => rgb <= "001000";
					when "011011101010101" => rgb <= "001000";
					when "011011101010110" => rgb <= "000000";
					when "011011101010111" => rgb <= "000000";
					when "011011101011000" => rgb <= "101111";
					when "011011101011001" => rgb <= "101111";
					when "011011101011010" => rgb <= "101111";
					when "011011101011011" => rgb <= "101111";
					when "011011101011100" => rgb <= "101111";
					when "011011101011101" => rgb <= "101111";
					when "011011101011110" => rgb <= "101111";
					when "011011101011111" => rgb <= "101111";
					when "011011101100000" => rgb <= "101111";
					when "011011101100001" => rgb <= "101111";
					when "011011101100010" => rgb <= "101111";
					when "011011101100011" => rgb <= "101111";
					when "011011101100100" => rgb <= "101111";
					when "011011101100101" => rgb <= "101111";
					when "011011101100110" => rgb <= "101111";
					when "011011101100111" => rgb <= "101111";
					when "011011101101000" => rgb <= "101111";
					when "011011101101001" => rgb <= "101111";
					when "011011101101010" => rgb <= "101111";
					when "011011101101011" => rgb <= "101111";
					when "011011101101100" => rgb <= "101111";
					when "011011101101101" => rgb <= "101111";
					when "011011101101110" => rgb <= "101111";
					when "011011101101111" => rgb <= "101111";
					when "011011101110000" => rgb <= "101111";
					when "011011101110001" => rgb <= "101111";
					when "011011101110010" => rgb <= "101111";
					when "011011101110011" => rgb <= "101111";
					when "011011101110100" => rgb <= "101111";
					when "011011101110101" => rgb <= "101111";
					when "011011101110110" => rgb <= "101111";
					when "011011101110111" => rgb <= "101111";
					when "011011101111000" => rgb <= "101111";
					when "011011101111001" => rgb <= "101111";
					when "011011101111010" => rgb <= "101111";
					when "011011101111011" => rgb <= "101111";
					when "011011101111100" => rgb <= "101111";
					when "011011101111101" => rgb <= "101111";
					when "011011101111110" => rgb <= "101111";
					when "011011101111111" => rgb <= "101111";
					when "011011110000000" => rgb <= "101111";
					when "011011110000001" => rgb <= "101111";
					when "011011110000010" => rgb <= "101111";
					when "011011110000011" => rgb <= "101111";
					when "011011110000100" => rgb <= "101111";
					when "011011110000101" => rgb <= "101111";
					when "011011110000110" => rgb <= "101111";
					when "011011110000111" => rgb <= "101111";
					when "011011110001000" => rgb <= "101111";
					when "011011110001001" => rgb <= "101111";
					when "011011110001010" => rgb <= "101111";
					when "011011110001011" => rgb <= "101111";
					when "011011110001100" => rgb <= "101111";
					when "011011110001101" => rgb <= "101111";
					when "011011110001110" => rgb <= "101111";
					when "011011110001111" => rgb <= "101111";
					when "011011110010000" => rgb <= "101111";
					when "011011110010001" => rgb <= "101111";
					when "011011110010010" => rgb <= "101111";
					when "011011110010011" => rgb <= "101111";
					when "011011110010100" => rgb <= "101111";
					when "011011110010101" => rgb <= "101111";
					when "011011110010110" => rgb <= "101111";
					when "011011110010111" => rgb <= "101111";
					when "011011110011000" => rgb <= "101111";
					when "011011110011001" => rgb <= "101111";
					when "011011110011010" => rgb <= "101111";
					when "011011110011011" => rgb <= "101111";
					when "011011110011100" => rgb <= "101111";
					when "011011110011101" => rgb <= "101111";
					when "011011110011110" => rgb <= "101111";
					when "011011110011111" => rgb <= "101111";
					when "011100000000000" => rgb <= "001000";
					when "011100000000001" => rgb <= "001000";
					when "011100000000010" => rgb <= "001000";
					when "011100000000011" => rgb <= "001000";
					when "011100000000100" => rgb <= "001000";
					when "011100000000101" => rgb <= "001000";
					when "011100000000110" => rgb <= "001000";
					when "011100000000111" => rgb <= "001000";
					when "011100000001000" => rgb <= "001000";
					when "011100000001001" => rgb <= "001000";
					when "011100000001010" => rgb <= "001000";
					when "011100000001011" => rgb <= "001000";
					when "011100000001100" => rgb <= "001000";
					when "011100000001101" => rgb <= "001000";
					when "011100000001110" => rgb <= "001000";
					when "011100000001111" => rgb <= "001000";
					when "011100000010000" => rgb <= "001000";
					when "011100000010001" => rgb <= "001000";
					when "011100000010010" => rgb <= "001000";
					when "011100000010011" => rgb <= "001000";
					when "011100000010100" => rgb <= "001000";
					when "011100000010101" => rgb <= "001000";
					when "011100000010110" => rgb <= "001000";
					when "011100000010111" => rgb <= "001000";
					when "011100000011000" => rgb <= "001000";
					when "011100000011001" => rgb <= "001000";
					when "011100000011010" => rgb <= "001000";
					when "011100000011011" => rgb <= "001000";
					when "011100000011100" => rgb <= "001000";
					when "011100000011101" => rgb <= "001000";
					when "011100000011110" => rgb <= "001000";
					when "011100000011111" => rgb <= "001000";
					when "011100000100000" => rgb <= "001000";
					when "011100000100001" => rgb <= "001000";
					when "011100000100010" => rgb <= "001000";
					when "011100000100011" => rgb <= "001000";
					when "011100000100100" => rgb <= "001000";
					when "011100000100101" => rgb <= "001000";
					when "011100000100110" => rgb <= "001000";
					when "011100000100111" => rgb <= "001000";
					when "011100000101000" => rgb <= "001000";
					when "011100000101001" => rgb <= "001000";
					when "011100000101010" => rgb <= "001000";
					when "011100000101011" => rgb <= "001000";
					when "011100000101100" => rgb <= "001000";
					when "011100000101101" => rgb <= "001000";
					when "011100000101110" => rgb <= "001000";
					when "011100000101111" => rgb <= "001000";
					when "011100000110000" => rgb <= "001000";
					when "011100000110001" => rgb <= "001000";
					when "011100000110010" => rgb <= "001000";
					when "011100000110011" => rgb <= "001000";
					when "011100000110100" => rgb <= "001000";
					when "011100000110101" => rgb <= "001000";
					when "011100000110110" => rgb <= "001000";
					when "011100000110111" => rgb <= "001000";
					when "011100000111000" => rgb <= "001000";
					when "011100000111001" => rgb <= "001000";
					when "011100000111010" => rgb <= "001000";
					when "011100000111011" => rgb <= "001000";
					when "011100000111100" => rgb <= "001000";
					when "011100000111101" => rgb <= "001000";
					when "011100000111110" => rgb <= "001000";
					when "011100000111111" => rgb <= "001000";
					when "011100001000000" => rgb <= "001000";
					when "011100001000001" => rgb <= "001000";
					when "011100001000010" => rgb <= "001000";
					when "011100001000011" => rgb <= "001000";
					when "011100001000100" => rgb <= "001000";
					when "011100001000101" => rgb <= "001000";
					when "011100001000110" => rgb <= "001000";
					when "011100001000111" => rgb <= "001000";
					when "011100001001000" => rgb <= "001000";
					when "011100001001001" => rgb <= "001000";
					when "011100001001010" => rgb <= "001000";
					when "011100001001011" => rgb <= "001000";
					when "011100001001100" => rgb <= "001000";
					when "011100001001101" => rgb <= "001000";
					when "011100001001110" => rgb <= "001000";
					when "011100001001111" => rgb <= "001000";
					when "011100001010000" => rgb <= "001000";
					when "011100001010001" => rgb <= "001000";
					when "011100001010010" => rgb <= "001000";
					when "011100001010011" => rgb <= "001000";
					when "011100001010100" => rgb <= "001000";
					when "011100001010101" => rgb <= "001000";
					when "011100001010110" => rgb <= "000000";
					when "011100001010111" => rgb <= "000000";
					when "011100001011000" => rgb <= "101111";
					when "011100001011001" => rgb <= "101111";
					when "011100001011010" => rgb <= "101111";
					when "011100001011011" => rgb <= "101111";
					when "011100001011100" => rgb <= "101111";
					when "011100001011101" => rgb <= "101111";
					when "011100001011110" => rgb <= "101111";
					when "011100001011111" => rgb <= "101111";
					when "011100001100000" => rgb <= "101111";
					when "011100001100001" => rgb <= "101111";
					when "011100001100010" => rgb <= "101111";
					when "011100001100011" => rgb <= "101111";
					when "011100001100100" => rgb <= "101111";
					when "011100001100101" => rgb <= "101111";
					when "011100001100110" => rgb <= "101111";
					when "011100001100111" => rgb <= "101111";
					when "011100001101000" => rgb <= "101111";
					when "011100001101001" => rgb <= "101111";
					when "011100001101010" => rgb <= "101111";
					when "011100001101011" => rgb <= "101111";
					when "011100001101100" => rgb <= "101111";
					when "011100001101101" => rgb <= "101111";
					when "011100001101110" => rgb <= "101111";
					when "011100001101111" => rgb <= "101111";
					when "011100001110000" => rgb <= "101111";
					when "011100001110001" => rgb <= "101111";
					when "011100001110010" => rgb <= "101111";
					when "011100001110011" => rgb <= "101111";
					when "011100001110100" => rgb <= "101111";
					when "011100001110101" => rgb <= "101111";
					when "011100001110110" => rgb <= "101111";
					when "011100001110111" => rgb <= "101111";
					when "011100001111000" => rgb <= "101111";
					when "011100001111001" => rgb <= "101111";
					when "011100001111010" => rgb <= "101111";
					when "011100001111011" => rgb <= "101111";
					when "011100001111100" => rgb <= "101111";
					when "011100001111101" => rgb <= "101111";
					when "011100001111110" => rgb <= "101111";
					when "011100001111111" => rgb <= "101111";
					when "011100010000000" => rgb <= "101111";
					when "011100010000001" => rgb <= "101111";
					when "011100010000010" => rgb <= "101111";
					when "011100010000011" => rgb <= "101111";
					when "011100010000100" => rgb <= "101111";
					when "011100010000101" => rgb <= "101111";
					when "011100010000110" => rgb <= "101111";
					when "011100010000111" => rgb <= "101111";
					when "011100010001000" => rgb <= "101111";
					when "011100010001001" => rgb <= "101111";
					when "011100010001010" => rgb <= "101111";
					when "011100010001011" => rgb <= "101111";
					when "011100010001100" => rgb <= "101111";
					when "011100010001101" => rgb <= "101111";
					when "011100010001110" => rgb <= "101111";
					when "011100010001111" => rgb <= "101111";
					when "011100010010000" => rgb <= "101111";
					when "011100010010001" => rgb <= "101111";
					when "011100010010010" => rgb <= "101111";
					when "011100010010011" => rgb <= "101111";
					when "011100010010100" => rgb <= "101111";
					when "011100010010101" => rgb <= "101111";
					when "011100010010110" => rgb <= "101111";
					when "011100010010111" => rgb <= "101111";
					when "011100010011000" => rgb <= "101111";
					when "011100010011001" => rgb <= "101111";
					when "011100010011010" => rgb <= "101111";
					when "011100010011011" => rgb <= "101111";
					when "011100010011100" => rgb <= "101111";
					when "011100010011101" => rgb <= "101111";
					when "011100010011110" => rgb <= "101111";
					when "011100010011111" => rgb <= "101111";
					when "011100100000000" => rgb <= "001000";
					when "011100100000001" => rgb <= "001000";
					when "011100100000010" => rgb <= "001000";
					when "011100100000011" => rgb <= "001000";
					when "011100100000100" => rgb <= "001000";
					when "011100100000101" => rgb <= "001000";
					when "011100100000110" => rgb <= "001000";
					when "011100100000111" => rgb <= "001000";
					when "011100100001000" => rgb <= "001000";
					when "011100100001001" => rgb <= "001000";
					when "011100100001010" => rgb <= "001000";
					when "011100100001011" => rgb <= "001000";
					when "011100100001100" => rgb <= "001000";
					when "011100100001101" => rgb <= "001000";
					when "011100100001110" => rgb <= "001000";
					when "011100100001111" => rgb <= "001000";
					when "011100100010000" => rgb <= "001000";
					when "011100100010001" => rgb <= "001000";
					when "011100100010010" => rgb <= "001000";
					when "011100100010011" => rgb <= "001000";
					when "011100100010100" => rgb <= "001000";
					when "011100100010101" => rgb <= "001000";
					when "011100100010110" => rgb <= "001000";
					when "011100100010111" => rgb <= "001000";
					when "011100100011000" => rgb <= "001000";
					when "011100100011001" => rgb <= "001000";
					when "011100100011010" => rgb <= "001000";
					when "011100100011011" => rgb <= "001000";
					when "011100100011100" => rgb <= "001000";
					when "011100100011101" => rgb <= "001000";
					when "011100100011110" => rgb <= "001000";
					when "011100100011111" => rgb <= "001000";
					when "011100100100000" => rgb <= "001000";
					when "011100100100001" => rgb <= "001000";
					when "011100100100010" => rgb <= "001000";
					when "011100100100011" => rgb <= "001000";
					when "011100100100100" => rgb <= "001000";
					when "011100100100101" => rgb <= "001000";
					when "011100100100110" => rgb <= "001000";
					when "011100100100111" => rgb <= "001000";
					when "011100100101000" => rgb <= "001000";
					when "011100100101001" => rgb <= "001000";
					when "011100100101010" => rgb <= "001000";
					when "011100100101011" => rgb <= "001000";
					when "011100100101100" => rgb <= "001000";
					when "011100100101101" => rgb <= "001000";
					when "011100100101110" => rgb <= "001000";
					when "011100100101111" => rgb <= "001000";
					when "011100100110000" => rgb <= "001000";
					when "011100100110001" => rgb <= "001000";
					when "011100100110010" => rgb <= "001000";
					when "011100100110011" => rgb <= "001000";
					when "011100100110100" => rgb <= "001000";
					when "011100100110101" => rgb <= "001000";
					when "011100100110110" => rgb <= "001000";
					when "011100100110111" => rgb <= "001000";
					when "011100100111000" => rgb <= "001000";
					when "011100100111001" => rgb <= "001000";
					when "011100100111010" => rgb <= "001000";
					when "011100100111011" => rgb <= "001000";
					when "011100100111100" => rgb <= "001000";
					when "011100100111101" => rgb <= "001000";
					when "011100100111110" => rgb <= "001000";
					when "011100100111111" => rgb <= "001000";
					when "011100101000000" => rgb <= "001000";
					when "011100101000001" => rgb <= "001000";
					when "011100101000010" => rgb <= "001000";
					when "011100101000011" => rgb <= "001000";
					when "011100101000100" => rgb <= "001000";
					when "011100101000101" => rgb <= "001000";
					when "011100101000110" => rgb <= "001000";
					when "011100101000111" => rgb <= "001000";
					when "011100101001000" => rgb <= "001000";
					when "011100101001001" => rgb <= "001000";
					when "011100101001010" => rgb <= "001000";
					when "011100101001011" => rgb <= "001000";
					when "011100101001100" => rgb <= "001000";
					when "011100101001101" => rgb <= "001000";
					when "011100101001110" => rgb <= "001000";
					when "011100101001111" => rgb <= "001000";
					when "011100101010000" => rgb <= "001000";
					when "011100101010001" => rgb <= "001000";
					when "011100101010010" => rgb <= "001000";
					when "011100101010011" => rgb <= "001000";
					when "011100101010100" => rgb <= "001000";
					when "011100101010101" => rgb <= "001000";
					when "011100101010110" => rgb <= "000000";
					when "011100101010111" => rgb <= "000000";
					when "011100101011000" => rgb <= "101111";
					when "011100101011001" => rgb <= "101111";
					when "011100101011010" => rgb <= "101111";
					when "011100101011011" => rgb <= "101111";
					when "011100101011100" => rgb <= "101111";
					when "011100101011101" => rgb <= "101111";
					when "011100101011110" => rgb <= "101111";
					when "011100101011111" => rgb <= "101111";
					when "011100101100000" => rgb <= "101111";
					when "011100101100001" => rgb <= "101111";
					when "011100101100010" => rgb <= "101111";
					when "011100101100011" => rgb <= "101111";
					when "011100101100100" => rgb <= "101111";
					when "011100101100101" => rgb <= "101111";
					when "011100101100110" => rgb <= "101111";
					when "011100101100111" => rgb <= "101111";
					when "011100101101000" => rgb <= "101111";
					when "011100101101001" => rgb <= "101111";
					when "011100101101010" => rgb <= "101111";
					when "011100101101011" => rgb <= "101111";
					when "011100101101100" => rgb <= "101111";
					when "011100101101101" => rgb <= "101111";
					when "011100101101110" => rgb <= "101111";
					when "011100101101111" => rgb <= "101111";
					when "011100101110000" => rgb <= "101111";
					when "011100101110001" => rgb <= "101111";
					when "011100101110010" => rgb <= "101111";
					when "011100101110011" => rgb <= "101111";
					when "011100101110100" => rgb <= "101111";
					when "011100101110101" => rgb <= "101111";
					when "011100101110110" => rgb <= "101111";
					when "011100101110111" => rgb <= "101111";
					when "011100101111000" => rgb <= "101111";
					when "011100101111001" => rgb <= "101111";
					when "011100101111010" => rgb <= "101111";
					when "011100101111011" => rgb <= "101111";
					when "011100101111100" => rgb <= "101111";
					when "011100101111101" => rgb <= "101111";
					when "011100101111110" => rgb <= "101111";
					when "011100101111111" => rgb <= "101111";
					when "011100110000000" => rgb <= "101111";
					when "011100110000001" => rgb <= "101111";
					when "011100110000010" => rgb <= "101111";
					when "011100110000011" => rgb <= "101111";
					when "011100110000100" => rgb <= "101111";
					when "011100110000101" => rgb <= "101111";
					when "011100110000110" => rgb <= "101111";
					when "011100110000111" => rgb <= "101111";
					when "011100110001000" => rgb <= "101111";
					when "011100110001001" => rgb <= "101111";
					when "011100110001010" => rgb <= "101111";
					when "011100110001011" => rgb <= "101111";
					when "011100110001100" => rgb <= "101111";
					when "011100110001101" => rgb <= "101111";
					when "011100110001110" => rgb <= "101111";
					when "011100110001111" => rgb <= "101111";
					when "011100110010000" => rgb <= "101111";
					when "011100110010001" => rgb <= "101111";
					when "011100110010010" => rgb <= "101111";
					when "011100110010011" => rgb <= "101111";
					when "011100110010100" => rgb <= "101111";
					when "011100110010101" => rgb <= "101111";
					when "011100110010110" => rgb <= "101111";
					when "011100110010111" => rgb <= "101111";
					when "011100110011000" => rgb <= "101111";
					when "011100110011001" => rgb <= "101111";
					when "011100110011010" => rgb <= "101111";
					when "011100110011011" => rgb <= "101111";
					when "011100110011100" => rgb <= "101111";
					when "011100110011101" => rgb <= "101111";
					when "011100110011110" => rgb <= "101111";
					when "011100110011111" => rgb <= "101111";
					when "011101000000000" => rgb <= "001000";
					when "011101000000001" => rgb <= "001000";
					when "011101000000010" => rgb <= "001000";
					when "011101000000011" => rgb <= "001000";
					when "011101000000100" => rgb <= "001000";
					when "011101000000101" => rgb <= "001000";
					when "011101000000110" => rgb <= "001000";
					when "011101000000111" => rgb <= "001000";
					when "011101000001000" => rgb <= "001000";
					when "011101000001001" => rgb <= "001000";
					when "011101000001010" => rgb <= "001000";
					when "011101000001011" => rgb <= "001000";
					when "011101000001100" => rgb <= "001000";
					when "011101000001101" => rgb <= "001000";
					when "011101000001110" => rgb <= "001000";
					when "011101000001111" => rgb <= "001000";
					when "011101000010000" => rgb <= "001000";
					when "011101000010001" => rgb <= "001000";
					when "011101000010010" => rgb <= "001000";
					when "011101000010011" => rgb <= "001000";
					when "011101000010100" => rgb <= "001000";
					when "011101000010101" => rgb <= "001000";
					when "011101000010110" => rgb <= "001000";
					when "011101000010111" => rgb <= "001000";
					when "011101000011000" => rgb <= "001000";
					when "011101000011001" => rgb <= "001000";
					when "011101000011010" => rgb <= "001000";
					when "011101000011011" => rgb <= "001000";
					when "011101000011100" => rgb <= "000000";
					when "011101000011101" => rgb <= "000000";
					when "011101000011110" => rgb <= "000000";
					when "011101000011111" => rgb <= "000000";
					when "011101000100000" => rgb <= "000000";
					when "011101000100001" => rgb <= "000000";
					when "011101000100010" => rgb <= "000000";
					when "011101000100011" => rgb <= "000000";
					when "011101000100100" => rgb <= "001000";
					when "011101000100101" => rgb <= "001000";
					when "011101000100110" => rgb <= "001000";
					when "011101000100111" => rgb <= "001000";
					when "011101000101000" => rgb <= "001000";
					when "011101000101001" => rgb <= "001000";
					when "011101000101010" => rgb <= "001000";
					when "011101000101011" => rgb <= "001000";
					when "011101000101100" => rgb <= "001000";
					when "011101000101101" => rgb <= "001000";
					when "011101000101110" => rgb <= "001000";
					when "011101000101111" => rgb <= "001000";
					when "011101000110000" => rgb <= "001000";
					when "011101000110001" => rgb <= "001000";
					when "011101000110010" => rgb <= "001000";
					when "011101000110011" => rgb <= "001000";
					when "011101000110100" => rgb <= "001000";
					when "011101000110101" => rgb <= "001000";
					when "011101000110110" => rgb <= "001000";
					when "011101000110111" => rgb <= "001000";
					when "011101000111000" => rgb <= "001000";
					when "011101000111001" => rgb <= "001000";
					when "011101000111010" => rgb <= "001000";
					when "011101000111011" => rgb <= "001000";
					when "011101000111100" => rgb <= "001000";
					when "011101000111101" => rgb <= "001000";
					when "011101000111110" => rgb <= "001000";
					when "011101000111111" => rgb <= "001000";
					when "011101001000000" => rgb <= "001000";
					when "011101001000001" => rgb <= "001000";
					when "011101001000010" => rgb <= "001000";
					when "011101001000011" => rgb <= "001000";
					when "011101001000100" => rgb <= "001000";
					when "011101001000101" => rgb <= "001000";
					when "011101001000110" => rgb <= "001000";
					when "011101001000111" => rgb <= "001000";
					when "011101001001000" => rgb <= "001000";
					when "011101001001001" => rgb <= "001000";
					when "011101001001010" => rgb <= "001000";
					when "011101001001011" => rgb <= "001000";
					when "011101001001100" => rgb <= "001000";
					when "011101001001101" => rgb <= "001000";
					when "011101001001110" => rgb <= "001000";
					when "011101001001111" => rgb <= "001000";
					when "011101001010000" => rgb <= "001000";
					when "011101001010001" => rgb <= "001000";
					when "011101001010010" => rgb <= "000000";
					when "011101001010011" => rgb <= "000000";
					when "011101001010100" => rgb <= "000000";
					when "011101001010101" => rgb <= "000000";
					when "011101001010110" => rgb <= "101111";
					when "011101001010111" => rgb <= "101111";
					when "011101001011000" => rgb <= "101111";
					when "011101001011001" => rgb <= "101111";
					when "011101001011010" => rgb <= "101111";
					when "011101001011011" => rgb <= "101111";
					when "011101001011100" => rgb <= "101111";
					when "011101001011101" => rgb <= "101111";
					when "011101001011110" => rgb <= "101111";
					when "011101001011111" => rgb <= "101111";
					when "011101001100000" => rgb <= "101111";
					when "011101001100001" => rgb <= "101111";
					when "011101001100010" => rgb <= "101111";
					when "011101001100011" => rgb <= "101111";
					when "011101001100100" => rgb <= "101111";
					when "011101001100101" => rgb <= "101111";
					when "011101001100110" => rgb <= "101111";
					when "011101001100111" => rgb <= "101111";
					when "011101001101000" => rgb <= "101111";
					when "011101001101001" => rgb <= "101111";
					when "011101001101010" => rgb <= "101111";
					when "011101001101011" => rgb <= "101111";
					when "011101001101100" => rgb <= "101111";
					when "011101001101101" => rgb <= "101111";
					when "011101001101110" => rgb <= "101111";
					when "011101001101111" => rgb <= "101111";
					when "011101001110000" => rgb <= "101111";
					when "011101001110001" => rgb <= "101111";
					when "011101001110010" => rgb <= "101111";
					when "011101001110011" => rgb <= "101111";
					when "011101001110100" => rgb <= "101111";
					when "011101001110101" => rgb <= "101111";
					when "011101001110110" => rgb <= "101111";
					when "011101001110111" => rgb <= "101111";
					when "011101001111000" => rgb <= "101111";
					when "011101001111001" => rgb <= "101111";
					when "011101001111010" => rgb <= "101111";
					when "011101001111011" => rgb <= "101111";
					when "011101001111100" => rgb <= "101111";
					when "011101001111101" => rgb <= "101111";
					when "011101001111110" => rgb <= "101111";
					when "011101001111111" => rgb <= "101111";
					when "011101010000000" => rgb <= "101111";
					when "011101010000001" => rgb <= "101111";
					when "011101010000010" => rgb <= "101111";
					when "011101010000011" => rgb <= "101111";
					when "011101010000100" => rgb <= "101111";
					when "011101010000101" => rgb <= "101111";
					when "011101010000110" => rgb <= "101111";
					when "011101010000111" => rgb <= "101111";
					when "011101010001000" => rgb <= "101111";
					when "011101010001001" => rgb <= "101111";
					when "011101010001010" => rgb <= "101111";
					when "011101010001011" => rgb <= "101111";
					when "011101010001100" => rgb <= "101111";
					when "011101010001101" => rgb <= "101111";
					when "011101010001110" => rgb <= "101111";
					when "011101010001111" => rgb <= "101111";
					when "011101010010000" => rgb <= "101111";
					when "011101010010001" => rgb <= "101111";
					when "011101010010010" => rgb <= "101111";
					when "011101010010011" => rgb <= "101111";
					when "011101010010100" => rgb <= "101111";
					when "011101010010101" => rgb <= "101111";
					when "011101010010110" => rgb <= "101111";
					when "011101010010111" => rgb <= "101111";
					when "011101010011000" => rgb <= "101111";
					when "011101010011001" => rgb <= "101111";
					when "011101010011010" => rgb <= "101111";
					when "011101010011011" => rgb <= "101111";
					when "011101010011100" => rgb <= "101111";
					when "011101010011101" => rgb <= "101111";
					when "011101010011110" => rgb <= "101111";
					when "011101010011111" => rgb <= "101111";
					when "011101100000000" => rgb <= "001000";
					when "011101100000001" => rgb <= "001000";
					when "011101100000010" => rgb <= "001000";
					when "011101100000011" => rgb <= "001000";
					when "011101100000100" => rgb <= "001000";
					when "011101100000101" => rgb <= "001000";
					when "011101100000110" => rgb <= "001000";
					when "011101100000111" => rgb <= "001000";
					when "011101100001000" => rgb <= "001000";
					when "011101100001001" => rgb <= "001000";
					when "011101100001010" => rgb <= "001000";
					when "011101100001011" => rgb <= "001000";
					when "011101100001100" => rgb <= "001000";
					when "011101100001101" => rgb <= "001000";
					when "011101100001110" => rgb <= "001000";
					when "011101100001111" => rgb <= "001000";
					when "011101100010000" => rgb <= "001000";
					when "011101100010001" => rgb <= "001000";
					when "011101100010010" => rgb <= "001000";
					when "011101100010011" => rgb <= "001000";
					when "011101100010100" => rgb <= "001000";
					when "011101100010101" => rgb <= "001000";
					when "011101100010110" => rgb <= "001000";
					when "011101100010111" => rgb <= "001000";
					when "011101100011000" => rgb <= "001000";
					when "011101100011001" => rgb <= "001000";
					when "011101100011010" => rgb <= "001000";
					when "011101100011011" => rgb <= "001000";
					when "011101100011100" => rgb <= "000000";
					when "011101100011101" => rgb <= "000000";
					when "011101100011110" => rgb <= "000000";
					when "011101100011111" => rgb <= "000000";
					when "011101100100000" => rgb <= "000000";
					when "011101100100001" => rgb <= "000000";
					when "011101100100010" => rgb <= "000000";
					when "011101100100011" => rgb <= "000000";
					when "011101100100100" => rgb <= "001000";
					when "011101100100101" => rgb <= "001000";
					when "011101100100110" => rgb <= "001000";
					when "011101100100111" => rgb <= "001000";
					when "011101100101000" => rgb <= "001000";
					when "011101100101001" => rgb <= "001000";
					when "011101100101010" => rgb <= "001000";
					when "011101100101011" => rgb <= "001000";
					when "011101100101100" => rgb <= "001000";
					when "011101100101101" => rgb <= "001000";
					when "011101100101110" => rgb <= "001000";
					when "011101100101111" => rgb <= "001000";
					when "011101100110000" => rgb <= "001000";
					when "011101100110001" => rgb <= "001000";
					when "011101100110010" => rgb <= "001000";
					when "011101100110011" => rgb <= "001000";
					when "011101100110100" => rgb <= "001000";
					when "011101100110101" => rgb <= "001000";
					when "011101100110110" => rgb <= "001000";
					when "011101100110111" => rgb <= "001000";
					when "011101100111000" => rgb <= "001000";
					when "011101100111001" => rgb <= "001000";
					when "011101100111010" => rgb <= "001000";
					when "011101100111011" => rgb <= "001000";
					when "011101100111100" => rgb <= "001000";
					when "011101100111101" => rgb <= "001000";
					when "011101100111110" => rgb <= "001000";
					when "011101100111111" => rgb <= "001000";
					when "011101101000000" => rgb <= "001000";
					when "011101101000001" => rgb <= "001000";
					when "011101101000010" => rgb <= "001000";
					when "011101101000011" => rgb <= "001000";
					when "011101101000100" => rgb <= "001000";
					when "011101101000101" => rgb <= "001000";
					when "011101101000110" => rgb <= "001000";
					when "011101101000111" => rgb <= "001000";
					when "011101101001000" => rgb <= "001000";
					when "011101101001001" => rgb <= "001000";
					when "011101101001010" => rgb <= "001000";
					when "011101101001011" => rgb <= "001000";
					when "011101101001100" => rgb <= "001000";
					when "011101101001101" => rgb <= "001000";
					when "011101101001110" => rgb <= "001000";
					when "011101101001111" => rgb <= "001000";
					when "011101101010000" => rgb <= "001000";
					when "011101101010001" => rgb <= "001000";
					when "011101101010010" => rgb <= "000000";
					when "011101101010011" => rgb <= "000000";
					when "011101101010100" => rgb <= "000000";
					when "011101101010101" => rgb <= "000000";
					when "011101101010110" => rgb <= "101111";
					when "011101101010111" => rgb <= "101111";
					when "011101101011000" => rgb <= "101111";
					when "011101101011001" => rgb <= "101111";
					when "011101101011010" => rgb <= "101111";
					when "011101101011011" => rgb <= "101111";
					when "011101101011100" => rgb <= "101111";
					when "011101101011101" => rgb <= "101111";
					when "011101101011110" => rgb <= "101111";
					when "011101101011111" => rgb <= "101111";
					when "011101101100000" => rgb <= "101111";
					when "011101101100001" => rgb <= "101111";
					when "011101101100010" => rgb <= "101111";
					when "011101101100011" => rgb <= "101111";
					when "011101101100100" => rgb <= "101111";
					when "011101101100101" => rgb <= "101111";
					when "011101101100110" => rgb <= "101111";
					when "011101101100111" => rgb <= "101111";
					when "011101101101000" => rgb <= "101111";
					when "011101101101001" => rgb <= "101111";
					when "011101101101010" => rgb <= "101111";
					when "011101101101011" => rgb <= "101111";
					when "011101101101100" => rgb <= "101111";
					when "011101101101101" => rgb <= "101111";
					when "011101101101110" => rgb <= "101111";
					when "011101101101111" => rgb <= "101111";
					when "011101101110000" => rgb <= "101111";
					when "011101101110001" => rgb <= "101111";
					when "011101101110010" => rgb <= "101111";
					when "011101101110011" => rgb <= "101111";
					when "011101101110100" => rgb <= "101111";
					when "011101101110101" => rgb <= "101111";
					when "011101101110110" => rgb <= "101111";
					when "011101101110111" => rgb <= "101111";
					when "011101101111000" => rgb <= "101111";
					when "011101101111001" => rgb <= "101111";
					when "011101101111010" => rgb <= "101111";
					when "011101101111011" => rgb <= "101111";
					when "011101101111100" => rgb <= "101111";
					when "011101101111101" => rgb <= "101111";
					when "011101101111110" => rgb <= "101111";
					when "011101101111111" => rgb <= "101111";
					when "011101110000000" => rgb <= "101111";
					when "011101110000001" => rgb <= "101111";
					when "011101110000010" => rgb <= "101111";
					when "011101110000011" => rgb <= "101111";
					when "011101110000100" => rgb <= "101111";
					when "011101110000101" => rgb <= "101111";
					when "011101110000110" => rgb <= "101111";
					when "011101110000111" => rgb <= "101111";
					when "011101110001000" => rgb <= "101111";
					when "011101110001001" => rgb <= "101111";
					when "011101110001010" => rgb <= "101111";
					when "011101110001011" => rgb <= "101111";
					when "011101110001100" => rgb <= "101111";
					when "011101110001101" => rgb <= "101111";
					when "011101110001110" => rgb <= "101111";
					when "011101110001111" => rgb <= "101111";
					when "011101110010000" => rgb <= "101111";
					when "011101110010001" => rgb <= "101111";
					when "011101110010010" => rgb <= "101111";
					when "011101110010011" => rgb <= "101111";
					when "011101110010100" => rgb <= "101111";
					when "011101110010101" => rgb <= "101111";
					when "011101110010110" => rgb <= "101111";
					when "011101110010111" => rgb <= "101111";
					when "011101110011000" => rgb <= "101111";
					when "011101110011001" => rgb <= "101111";
					when "011101110011010" => rgb <= "101111";
					when "011101110011011" => rgb <= "101111";
					when "011101110011100" => rgb <= "101111";
					when "011101110011101" => rgb <= "101111";
					when "011101110011110" => rgb <= "101111";
					when "011101110011111" => rgb <= "101111";
					when "011110000000000" => rgb <= "001000";
					when "011110000000001" => rgb <= "001000";
					when "011110000000010" => rgb <= "001000";
					when "011110000000011" => rgb <= "001000";
					when "011110000000100" => rgb <= "001000";
					when "011110000000101" => rgb <= "001000";
					when "011110000000110" => rgb <= "001000";
					when "011110000000111" => rgb <= "001000";
					when "011110000001000" => rgb <= "001000";
					when "011110000001001" => rgb <= "001000";
					when "011110000001010" => rgb <= "001000";
					when "011110000001011" => rgb <= "001000";
					when "011110000001100" => rgb <= "001000";
					when "011110000001101" => rgb <= "001000";
					when "011110000001110" => rgb <= "001000";
					when "011110000001111" => rgb <= "001000";
					when "011110000010000" => rgb <= "001000";
					when "011110000010001" => rgb <= "001000";
					when "011110000010010" => rgb <= "001000";
					when "011110000010011" => rgb <= "001000";
					when "011110000010100" => rgb <= "001000";
					when "011110000010101" => rgb <= "001000";
					when "011110000010110" => rgb <= "001000";
					when "011110000010111" => rgb <= "001000";
					when "011110000011000" => rgb <= "001000";
					when "011110000011001" => rgb <= "001000";
					when "011110000011010" => rgb <= "000000";
					when "011110000011011" => rgb <= "000000";
					when "011110000011100" => rgb <= "000000";
					when "011110000011101" => rgb <= "000000";
					when "011110000011110" => rgb <= "101111";
					when "011110000011111" => rgb <= "101111";
					when "011110000100000" => rgb <= "000000";
					when "011110000100001" => rgb <= "000000";
					when "011110000100010" => rgb <= "010000";
					when "011110000100011" => rgb <= "010000";
					when "011110000100100" => rgb <= "000000";
					when "011110000100101" => rgb <= "000000";
					when "011110000100110" => rgb <= "000000";
					when "011110000100111" => rgb <= "000000";
					when "011110000101000" => rgb <= "001000";
					when "011110000101001" => rgb <= "001000";
					when "011110000101010" => rgb <= "001000";
					when "011110000101011" => rgb <= "001000";
					when "011110000101100" => rgb <= "000000";
					when "011110000101101" => rgb <= "000000";
					when "011110000101110" => rgb <= "000000";
					when "011110000101111" => rgb <= "000000";
					when "011110000110000" => rgb <= "001000";
					when "011110000110001" => rgb <= "001000";
					when "011110000110010" => rgb <= "000000";
					when "011110000110011" => rgb <= "000000";
					when "011110000110100" => rgb <= "000000";
					when "011110000110101" => rgb <= "000000";
					when "011110000110110" => rgb <= "000000";
					when "011110000110111" => rgb <= "000000";
					when "011110000111000" => rgb <= "001000";
					when "011110000111001" => rgb <= "001000";
					when "011110000111010" => rgb <= "001000";
					when "011110000111011" => rgb <= "001000";
					when "011110000111100" => rgb <= "001000";
					when "011110000111101" => rgb <= "001000";
					when "011110000111110" => rgb <= "001000";
					when "011110000111111" => rgb <= "001000";
					when "011110001000000" => rgb <= "001000";
					when "011110001000001" => rgb <= "001000";
					when "011110001000010" => rgb <= "001000";
					when "011110001000011" => rgb <= "001000";
					when "011110001000100" => rgb <= "001000";
					when "011110001000101" => rgb <= "001000";
					when "011110001000110" => rgb <= "001000";
					when "011110001000111" => rgb <= "001000";
					when "011110001001000" => rgb <= "001000";
					when "011110001001001" => rgb <= "001000";
					when "011110001001010" => rgb <= "001000";
					when "011110001001011" => rgb <= "001000";
					when "011110001001100" => rgb <= "001000";
					when "011110001001101" => rgb <= "001000";
					when "011110001001110" => rgb <= "001000";
					when "011110001001111" => rgb <= "001000";
					when "011110001010000" => rgb <= "000000";
					when "011110001010001" => rgb <= "000000";
					when "011110001010010" => rgb <= "000000";
					when "011110001010011" => rgb <= "000000";
					when "011110001010100" => rgb <= "101111";
					when "011110001010101" => rgb <= "101111";
					when "011110001010110" => rgb <= "101111";
					when "011110001010111" => rgb <= "101111";
					when "011110001011000" => rgb <= "101111";
					when "011110001011001" => rgb <= "101111";
					when "011110001011010" => rgb <= "101111";
					when "011110001011011" => rgb <= "101111";
					when "011110001011100" => rgb <= "101111";
					when "011110001011101" => rgb <= "101111";
					when "011110001011110" => rgb <= "101111";
					when "011110001011111" => rgb <= "101111";
					when "011110001100000" => rgb <= "101111";
					when "011110001100001" => rgb <= "101111";
					when "011110001100010" => rgb <= "101111";
					when "011110001100011" => rgb <= "101111";
					when "011110001100100" => rgb <= "101111";
					when "011110001100101" => rgb <= "101111";
					when "011110001100110" => rgb <= "101111";
					when "011110001100111" => rgb <= "101111";
					when "011110001101000" => rgb <= "101111";
					when "011110001101001" => rgb <= "101111";
					when "011110001101010" => rgb <= "101111";
					when "011110001101011" => rgb <= "101111";
					when "011110001101100" => rgb <= "101111";
					when "011110001101101" => rgb <= "101111";
					when "011110001101110" => rgb <= "101111";
					when "011110001101111" => rgb <= "101111";
					when "011110001110000" => rgb <= "101111";
					when "011110001110001" => rgb <= "101111";
					when "011110001110010" => rgb <= "101111";
					when "011110001110011" => rgb <= "101111";
					when "011110001110100" => rgb <= "101111";
					when "011110001110101" => rgb <= "101111";
					when "011110001110110" => rgb <= "101111";
					when "011110001110111" => rgb <= "101111";
					when "011110001111000" => rgb <= "101111";
					when "011110001111001" => rgb <= "101111";
					when "011110001111010" => rgb <= "101111";
					when "011110001111011" => rgb <= "101111";
					when "011110001111100" => rgb <= "101111";
					when "011110001111101" => rgb <= "101111";
					when "011110001111110" => rgb <= "101111";
					when "011110001111111" => rgb <= "101111";
					when "011110010000000" => rgb <= "101111";
					when "011110010000001" => rgb <= "101111";
					when "011110010000010" => rgb <= "101111";
					when "011110010000011" => rgb <= "101111";
					when "011110010000100" => rgb <= "101111";
					when "011110010000101" => rgb <= "101111";
					when "011110010000110" => rgb <= "101111";
					when "011110010000111" => rgb <= "101111";
					when "011110010001000" => rgb <= "101111";
					when "011110010001001" => rgb <= "101111";
					when "011110010001010" => rgb <= "101111";
					when "011110010001011" => rgb <= "101111";
					when "011110010001100" => rgb <= "101111";
					when "011110010001101" => rgb <= "101111";
					when "011110010001110" => rgb <= "101111";
					when "011110010001111" => rgb <= "101111";
					when "011110010010000" => rgb <= "101111";
					when "011110010010001" => rgb <= "101111";
					when "011110010010010" => rgb <= "101111";
					when "011110010010011" => rgb <= "101111";
					when "011110010010100" => rgb <= "101111";
					when "011110010010101" => rgb <= "101111";
					when "011110010010110" => rgb <= "101111";
					when "011110010010111" => rgb <= "101111";
					when "011110010011000" => rgb <= "101111";
					when "011110010011001" => rgb <= "101111";
					when "011110010011010" => rgb <= "101111";
					when "011110010011011" => rgb <= "101111";
					when "011110010011100" => rgb <= "101111";
					when "011110010011101" => rgb <= "101111";
					when "011110010011110" => rgb <= "101111";
					when "011110010011111" => rgb <= "101111";
					when "011110100000000" => rgb <= "001000";
					when "011110100000001" => rgb <= "001000";
					when "011110100000010" => rgb <= "001000";
					when "011110100000011" => rgb <= "001000";
					when "011110100000100" => rgb <= "001000";
					when "011110100000101" => rgb <= "001000";
					when "011110100000110" => rgb <= "001000";
					when "011110100000111" => rgb <= "001000";
					when "011110100001000" => rgb <= "001000";
					when "011110100001001" => rgb <= "001000";
					when "011110100001010" => rgb <= "001000";
					when "011110100001011" => rgb <= "001000";
					when "011110100001100" => rgb <= "001000";
					when "011110100001101" => rgb <= "001000";
					when "011110100001110" => rgb <= "001000";
					when "011110100001111" => rgb <= "001000";
					when "011110100010000" => rgb <= "001000";
					when "011110100010001" => rgb <= "001000";
					when "011110100010010" => rgb <= "001000";
					when "011110100010011" => rgb <= "001000";
					when "011110100010100" => rgb <= "001000";
					when "011110100010101" => rgb <= "001000";
					when "011110100010110" => rgb <= "001000";
					when "011110100010111" => rgb <= "001000";
					when "011110100011000" => rgb <= "001000";
					when "011110100011001" => rgb <= "001000";
					when "011110100011010" => rgb <= "000000";
					when "011110100011011" => rgb <= "000000";
					when "011110100011100" => rgb <= "000000";
					when "011110100011101" => rgb <= "000000";
					when "011110100011110" => rgb <= "101111";
					when "011110100011111" => rgb <= "101111";
					when "011110100100000" => rgb <= "000000";
					when "011110100100001" => rgb <= "000000";
					when "011110100100010" => rgb <= "010000";
					when "011110100100011" => rgb <= "010000";
					when "011110100100100" => rgb <= "000000";
					when "011110100100101" => rgb <= "000000";
					when "011110100100110" => rgb <= "000000";
					when "011110100100111" => rgb <= "000000";
					when "011110100101000" => rgb <= "001000";
					when "011110100101001" => rgb <= "001000";
					when "011110100101010" => rgb <= "001000";
					when "011110100101011" => rgb <= "001000";
					when "011110100101100" => rgb <= "000000";
					when "011110100101101" => rgb <= "000000";
					when "011110100101110" => rgb <= "000000";
					when "011110100101111" => rgb <= "000000";
					when "011110100110000" => rgb <= "001000";
					when "011110100110001" => rgb <= "001000";
					when "011110100110010" => rgb <= "000000";
					when "011110100110011" => rgb <= "000000";
					when "011110100110100" => rgb <= "000000";
					when "011110100110101" => rgb <= "000000";
					when "011110100110110" => rgb <= "000000";
					when "011110100110111" => rgb <= "000000";
					when "011110100111000" => rgb <= "001000";
					when "011110100111001" => rgb <= "001000";
					when "011110100111010" => rgb <= "001000";
					when "011110100111011" => rgb <= "001000";
					when "011110100111100" => rgb <= "001000";
					when "011110100111101" => rgb <= "001000";
					when "011110100111110" => rgb <= "001000";
					when "011110100111111" => rgb <= "001000";
					when "011110101000000" => rgb <= "001000";
					when "011110101000001" => rgb <= "001000";
					when "011110101000010" => rgb <= "001000";
					when "011110101000011" => rgb <= "001000";
					when "011110101000100" => rgb <= "001000";
					when "011110101000101" => rgb <= "001000";
					when "011110101000110" => rgb <= "001000";
					when "011110101000111" => rgb <= "001000";
					when "011110101001000" => rgb <= "001000";
					when "011110101001001" => rgb <= "001000";
					when "011110101001010" => rgb <= "001000";
					when "011110101001011" => rgb <= "001000";
					when "011110101001100" => rgb <= "001000";
					when "011110101001101" => rgb <= "001000";
					when "011110101001110" => rgb <= "001000";
					when "011110101001111" => rgb <= "001000";
					when "011110101010000" => rgb <= "000000";
					when "011110101010001" => rgb <= "000000";
					when "011110101010010" => rgb <= "000000";
					when "011110101010011" => rgb <= "000000";
					when "011110101010100" => rgb <= "101111";
					when "011110101010101" => rgb <= "101111";
					when "011110101010110" => rgb <= "101111";
					when "011110101010111" => rgb <= "101111";
					when "011110101011000" => rgb <= "101111";
					when "011110101011001" => rgb <= "101111";
					when "011110101011010" => rgb <= "101111";
					when "011110101011011" => rgb <= "101111";
					when "011110101011100" => rgb <= "101111";
					when "011110101011101" => rgb <= "101111";
					when "011110101011110" => rgb <= "101111";
					when "011110101011111" => rgb <= "101111";
					when "011110101100000" => rgb <= "101111";
					when "011110101100001" => rgb <= "101111";
					when "011110101100010" => rgb <= "101111";
					when "011110101100011" => rgb <= "101111";
					when "011110101100100" => rgb <= "101111";
					when "011110101100101" => rgb <= "101111";
					when "011110101100110" => rgb <= "101111";
					when "011110101100111" => rgb <= "101111";
					when "011110101101000" => rgb <= "101111";
					when "011110101101001" => rgb <= "101111";
					when "011110101101010" => rgb <= "101111";
					when "011110101101011" => rgb <= "101111";
					when "011110101101100" => rgb <= "101111";
					when "011110101101101" => rgb <= "101111";
					when "011110101101110" => rgb <= "101111";
					when "011110101101111" => rgb <= "101111";
					when "011110101110000" => rgb <= "101111";
					when "011110101110001" => rgb <= "101111";
					when "011110101110010" => rgb <= "101111";
					when "011110101110011" => rgb <= "101111";
					when "011110101110100" => rgb <= "101111";
					when "011110101110101" => rgb <= "101111";
					when "011110101110110" => rgb <= "101111";
					when "011110101110111" => rgb <= "101111";
					when "011110101111000" => rgb <= "101111";
					when "011110101111001" => rgb <= "101111";
					when "011110101111010" => rgb <= "101111";
					when "011110101111011" => rgb <= "101111";
					when "011110101111100" => rgb <= "101111";
					when "011110101111101" => rgb <= "101111";
					when "011110101111110" => rgb <= "101111";
					when "011110101111111" => rgb <= "101111";
					when "011110110000000" => rgb <= "101111";
					when "011110110000001" => rgb <= "101111";
					when "011110110000010" => rgb <= "101111";
					when "011110110000011" => rgb <= "101111";
					when "011110110000100" => rgb <= "101111";
					when "011110110000101" => rgb <= "101111";
					when "011110110000110" => rgb <= "101111";
					when "011110110000111" => rgb <= "101111";
					when "011110110001000" => rgb <= "101111";
					when "011110110001001" => rgb <= "101111";
					when "011110110001010" => rgb <= "101111";
					when "011110110001011" => rgb <= "101111";
					when "011110110001100" => rgb <= "101111";
					when "011110110001101" => rgb <= "101111";
					when "011110110001110" => rgb <= "101111";
					when "011110110001111" => rgb <= "101111";
					when "011110110010000" => rgb <= "101111";
					when "011110110010001" => rgb <= "101111";
					when "011110110010010" => rgb <= "101111";
					when "011110110010011" => rgb <= "101111";
					when "011110110010100" => rgb <= "101111";
					when "011110110010101" => rgb <= "101111";
					when "011110110010110" => rgb <= "101111";
					when "011110110010111" => rgb <= "101111";
					when "011110110011000" => rgb <= "101111";
					when "011110110011001" => rgb <= "101111";
					when "011110110011010" => rgb <= "101111";
					when "011110110011011" => rgb <= "101111";
					when "011110110011100" => rgb <= "101111";
					when "011110110011101" => rgb <= "101111";
					when "011110110011110" => rgb <= "101111";
					when "011110110011111" => rgb <= "101111";
					when "011111000000000" => rgb <= "001000";
					when "011111000000001" => rgb <= "001000";
					when "011111000000010" => rgb <= "001000";
					when "011111000000011" => rgb <= "001000";
					when "011111000000100" => rgb <= "001000";
					when "011111000000101" => rgb <= "001000";
					when "011111000000110" => rgb <= "001000";
					when "011111000000111" => rgb <= "001000";
					when "011111000001000" => rgb <= "000000";
					when "011111000001001" => rgb <= "000000";
					when "011111000001010" => rgb <= "000000";
					when "011111000001011" => rgb <= "000000";
					when "011111000001100" => rgb <= "000000";
					when "011111000001101" => rgb <= "000000";
					when "011111000001110" => rgb <= "001000";
					when "011111000001111" => rgb <= "001000";
					when "011111000010000" => rgb <= "001000";
					when "011111000010001" => rgb <= "001000";
					when "011111000010010" => rgb <= "001000";
					when "011111000010011" => rgb <= "001000";
					when "011111000010100" => rgb <= "000000";
					when "011111000010101" => rgb <= "000000";
					when "011111000010110" => rgb <= "000000";
					when "011111000010111" => rgb <= "000000";
					when "011111000011000" => rgb <= "000000";
					when "011111000011001" => rgb <= "000000";
					when "011111000011010" => rgb <= "101111";
					when "011111000011011" => rgb <= "101111";
					when "011111000011100" => rgb <= "101111";
					when "011111000011101" => rgb <= "101111";
					when "011111000011110" => rgb <= "101111";
					when "011111000011111" => rgb <= "101111";
					when "011111000100000" => rgb <= "000000";
					when "011111000100001" => rgb <= "000000";
					when "011111000100010" => rgb <= "010000";
					when "011111000100011" => rgb <= "010000";
					when "011111000100100" => rgb <= "010000";
					when "011111000100101" => rgb <= "010000";
					when "011111000100110" => rgb <= "000000";
					when "011111000100111" => rgb <= "000000";
					when "011111000101000" => rgb <= "000000";
					when "011111000101001" => rgb <= "000000";
					when "011111000101010" => rgb <= "000000";
					when "011111000101011" => rgb <= "000000";
					when "011111000101100" => rgb <= "010000";
					when "011111000101101" => rgb <= "010000";
					when "011111000101110" => rgb <= "010000";
					when "011111000101111" => rgb <= "010000";
					when "011111000110000" => rgb <= "000000";
					when "011111000110001" => rgb <= "000000";
					when "011111000110010" => rgb <= "010000";
					when "011111000110011" => rgb <= "010000";
					when "011111000110100" => rgb <= "000000";
					when "011111000110101" => rgb <= "000000";
					when "011111000110110" => rgb <= "101111";
					when "011111000110111" => rgb <= "101111";
					when "011111000111000" => rgb <= "000000";
					when "011111000111001" => rgb <= "000000";
					when "011111000111010" => rgb <= "000000";
					when "011111000111011" => rgb <= "000000";
					when "011111000111100" => rgb <= "000000";
					when "011111000111101" => rgb <= "000000";
					when "011111000111110" => rgb <= "001000";
					when "011111000111111" => rgb <= "001000";
					when "011111001000000" => rgb <= "001000";
					when "011111001000001" => rgb <= "001000";
					when "011111001000010" => rgb <= "001000";
					when "011111001000011" => rgb <= "001000";
					when "011111001000100" => rgb <= "001000";
					when "011111001000101" => rgb <= "001000";
					when "011111001000110" => rgb <= "001000";
					when "011111001000111" => rgb <= "001000";
					when "011111001001000" => rgb <= "001000";
					when "011111001001001" => rgb <= "001000";
					when "011111001001010" => rgb <= "001000";
					when "011111001001011" => rgb <= "001000";
					when "011111001001100" => rgb <= "001000";
					when "011111001001101" => rgb <= "001000";
					when "011111001001110" => rgb <= "000000";
					when "011111001001111" => rgb <= "000000";
					when "011111001010000" => rgb <= "000000";
					when "011111001010001" => rgb <= "000000";
					when "011111001010010" => rgb <= "101111";
					when "011111001010011" => rgb <= "101111";
					when "011111001010100" => rgb <= "101111";
					when "011111001010101" => rgb <= "101111";
					when "011111001010110" => rgb <= "101111";
					when "011111001010111" => rgb <= "101111";
					when "011111001011000" => rgb <= "101111";
					when "011111001011001" => rgb <= "101111";
					when "011111001011010" => rgb <= "101111";
					when "011111001011011" => rgb <= "101111";
					when "011111001011100" => rgb <= "101111";
					when "011111001011101" => rgb <= "101111";
					when "011111001011110" => rgb <= "101111";
					when "011111001011111" => rgb <= "101111";
					when "011111001100000" => rgb <= "101111";
					when "011111001100001" => rgb <= "101111";
					when "011111001100010" => rgb <= "101111";
					when "011111001100011" => rgb <= "101111";
					when "011111001100100" => rgb <= "101111";
					when "011111001100101" => rgb <= "101111";
					when "011111001100110" => rgb <= "101111";
					when "011111001100111" => rgb <= "101111";
					when "011111001101000" => rgb <= "101111";
					when "011111001101001" => rgb <= "101111";
					when "011111001101010" => rgb <= "101111";
					when "011111001101011" => rgb <= "101111";
					when "011111001101100" => rgb <= "101111";
					when "011111001101101" => rgb <= "101111";
					when "011111001101110" => rgb <= "101111";
					when "011111001101111" => rgb <= "101111";
					when "011111001110000" => rgb <= "101111";
					when "011111001110001" => rgb <= "101111";
					when "011111001110010" => rgb <= "101111";
					when "011111001110011" => rgb <= "101111";
					when "011111001110100" => rgb <= "101111";
					when "011111001110101" => rgb <= "101111";
					when "011111001110110" => rgb <= "101111";
					when "011111001110111" => rgb <= "101111";
					when "011111001111000" => rgb <= "101111";
					when "011111001111001" => rgb <= "101111";
					when "011111001111010" => rgb <= "101111";
					when "011111001111011" => rgb <= "101111";
					when "011111001111100" => rgb <= "101111";
					when "011111001111101" => rgb <= "101111";
					when "011111001111110" => rgb <= "101111";
					when "011111001111111" => rgb <= "101111";
					when "011111010000000" => rgb <= "101111";
					when "011111010000001" => rgb <= "101111";
					when "011111010000010" => rgb <= "101111";
					when "011111010000011" => rgb <= "101111";
					when "011111010000100" => rgb <= "101111";
					when "011111010000101" => rgb <= "101111";
					when "011111010000110" => rgb <= "101111";
					when "011111010000111" => rgb <= "101111";
					when "011111010001000" => rgb <= "101111";
					when "011111010001001" => rgb <= "101111";
					when "011111010001010" => rgb <= "101111";
					when "011111010001011" => rgb <= "101111";
					when "011111010001100" => rgb <= "101111";
					when "011111010001101" => rgb <= "101111";
					when "011111010001110" => rgb <= "101111";
					when "011111010001111" => rgb <= "101111";
					when "011111010010000" => rgb <= "101111";
					when "011111010010001" => rgb <= "101111";
					when "011111010010010" => rgb <= "101111";
					when "011111010010011" => rgb <= "101111";
					when "011111010010100" => rgb <= "101111";
					when "011111010010101" => rgb <= "101111";
					when "011111010010110" => rgb <= "101111";
					when "011111010010111" => rgb <= "101111";
					when "011111010011000" => rgb <= "101111";
					when "011111010011001" => rgb <= "101111";
					when "011111010011010" => rgb <= "101111";
					when "011111010011011" => rgb <= "101111";
					when "011111010011100" => rgb <= "101111";
					when "011111010011101" => rgb <= "101111";
					when "011111010011110" => rgb <= "101111";
					when "011111010011111" => rgb <= "101111";
					when "011111100000000" => rgb <= "001000";
					when "011111100000001" => rgb <= "001000";
					when "011111100000010" => rgb <= "001000";
					when "011111100000011" => rgb <= "001000";
					when "011111100000100" => rgb <= "001000";
					when "011111100000101" => rgb <= "001000";
					when "011111100000110" => rgb <= "001000";
					when "011111100000111" => rgb <= "001000";
					when "011111100001000" => rgb <= "000000";
					when "011111100001001" => rgb <= "000000";
					when "011111100001010" => rgb <= "000000";
					when "011111100001011" => rgb <= "000000";
					when "011111100001100" => rgb <= "000000";
					when "011111100001101" => rgb <= "000000";
					when "011111100001110" => rgb <= "001000";
					when "011111100001111" => rgb <= "001000";
					when "011111100010000" => rgb <= "001000";
					when "011111100010001" => rgb <= "001000";
					when "011111100010010" => rgb <= "001000";
					when "011111100010011" => rgb <= "001000";
					when "011111100010100" => rgb <= "000000";
					when "011111100010101" => rgb <= "000000";
					when "011111100010110" => rgb <= "000000";
					when "011111100010111" => rgb <= "000000";
					when "011111100011000" => rgb <= "000000";
					when "011111100011001" => rgb <= "000000";
					when "011111100011010" => rgb <= "101111";
					when "011111100011011" => rgb <= "101111";
					when "011111100011100" => rgb <= "101111";
					when "011111100011101" => rgb <= "101111";
					when "011111100011110" => rgb <= "101111";
					when "011111100011111" => rgb <= "101111";
					when "011111100100000" => rgb <= "000000";
					when "011111100100001" => rgb <= "000000";
					when "011111100100010" => rgb <= "010000";
					when "011111100100011" => rgb <= "010000";
					when "011111100100100" => rgb <= "010000";
					when "011111100100101" => rgb <= "010000";
					when "011111100100110" => rgb <= "000000";
					when "011111100100111" => rgb <= "000000";
					when "011111100101000" => rgb <= "000000";
					when "011111100101001" => rgb <= "000000";
					when "011111100101010" => rgb <= "000000";
					when "011111100101011" => rgb <= "000000";
					when "011111100101100" => rgb <= "010000";
					when "011111100101101" => rgb <= "010000";
					when "011111100101110" => rgb <= "010000";
					when "011111100101111" => rgb <= "010000";
					when "011111100110000" => rgb <= "000000";
					when "011111100110001" => rgb <= "000000";
					when "011111100110010" => rgb <= "010000";
					when "011111100110011" => rgb <= "010000";
					when "011111100110100" => rgb <= "000000";
					when "011111100110101" => rgb <= "000000";
					when "011111100110110" => rgb <= "101111";
					when "011111100110111" => rgb <= "101111";
					when "011111100111000" => rgb <= "000000";
					when "011111100111001" => rgb <= "000000";
					when "011111100111010" => rgb <= "000000";
					when "011111100111011" => rgb <= "000000";
					when "011111100111100" => rgb <= "000000";
					when "011111100111101" => rgb <= "000000";
					when "011111100111110" => rgb <= "001000";
					when "011111100111111" => rgb <= "001000";
					when "011111101000000" => rgb <= "001000";
					when "011111101000001" => rgb <= "001000";
					when "011111101000010" => rgb <= "001000";
					when "011111101000011" => rgb <= "001000";
					when "011111101000100" => rgb <= "001000";
					when "011111101000101" => rgb <= "001000";
					when "011111101000110" => rgb <= "001000";
					when "011111101000111" => rgb <= "001000";
					when "011111101001000" => rgb <= "001000";
					when "011111101001001" => rgb <= "001000";
					when "011111101001010" => rgb <= "001000";
					when "011111101001011" => rgb <= "001000";
					when "011111101001100" => rgb <= "001000";
					when "011111101001101" => rgb <= "001000";
					when "011111101001110" => rgb <= "000000";
					when "011111101001111" => rgb <= "000000";
					when "011111101010000" => rgb <= "000000";
					when "011111101010001" => rgb <= "000000";
					when "011111101010010" => rgb <= "101111";
					when "011111101010011" => rgb <= "101111";
					when "011111101010100" => rgb <= "101111";
					when "011111101010101" => rgb <= "101111";
					when "011111101010110" => rgb <= "101111";
					when "011111101010111" => rgb <= "101111";
					when "011111101011000" => rgb <= "101111";
					when "011111101011001" => rgb <= "101111";
					when "011111101011010" => rgb <= "101111";
					when "011111101011011" => rgb <= "101111";
					when "011111101011100" => rgb <= "101111";
					when "011111101011101" => rgb <= "101111";
					when "011111101011110" => rgb <= "101111";
					when "011111101011111" => rgb <= "101111";
					when "011111101100000" => rgb <= "101111";
					when "011111101100001" => rgb <= "101111";
					when "011111101100010" => rgb <= "101111";
					when "011111101100011" => rgb <= "101111";
					when "011111101100100" => rgb <= "101111";
					when "011111101100101" => rgb <= "101111";
					when "011111101100110" => rgb <= "101111";
					when "011111101100111" => rgb <= "101111";
					when "011111101101000" => rgb <= "101111";
					when "011111101101001" => rgb <= "101111";
					when "011111101101010" => rgb <= "101111";
					when "011111101101011" => rgb <= "101111";
					when "011111101101100" => rgb <= "101111";
					when "011111101101101" => rgb <= "101111";
					when "011111101101110" => rgb <= "101111";
					when "011111101101111" => rgb <= "101111";
					when "011111101110000" => rgb <= "101111";
					when "011111101110001" => rgb <= "101111";
					when "011111101110010" => rgb <= "101111";
					when "011111101110011" => rgb <= "101111";
					when "011111101110100" => rgb <= "101111";
					when "011111101110101" => rgb <= "101111";
					when "011111101110110" => rgb <= "101111";
					when "011111101110111" => rgb <= "101111";
					when "011111101111000" => rgb <= "101111";
					when "011111101111001" => rgb <= "101111";
					when "011111101111010" => rgb <= "101111";
					when "011111101111011" => rgb <= "101111";
					when "011111101111100" => rgb <= "101111";
					when "011111101111101" => rgb <= "101111";
					when "011111101111110" => rgb <= "101111";
					when "011111101111111" => rgb <= "101111";
					when "011111110000000" => rgb <= "101111";
					when "011111110000001" => rgb <= "101111";
					when "011111110000010" => rgb <= "101111";
					when "011111110000011" => rgb <= "101111";
					when "011111110000100" => rgb <= "101111";
					when "011111110000101" => rgb <= "101111";
					when "011111110000110" => rgb <= "101111";
					when "011111110000111" => rgb <= "101111";
					when "011111110001000" => rgb <= "101111";
					when "011111110001001" => rgb <= "101111";
					when "011111110001010" => rgb <= "101111";
					when "011111110001011" => rgb <= "101111";
					when "011111110001100" => rgb <= "101111";
					when "011111110001101" => rgb <= "101111";
					when "011111110001110" => rgb <= "101111";
					when "011111110001111" => rgb <= "101111";
					when "011111110010000" => rgb <= "101111";
					when "011111110010001" => rgb <= "101111";
					when "011111110010010" => rgb <= "101111";
					when "011111110010011" => rgb <= "101111";
					when "011111110010100" => rgb <= "101111";
					when "011111110010101" => rgb <= "101111";
					when "011111110010110" => rgb <= "101111";
					when "011111110010111" => rgb <= "101111";
					when "011111110011000" => rgb <= "101111";
					when "011111110011001" => rgb <= "101111";
					when "011111110011010" => rgb <= "101111";
					when "011111110011011" => rgb <= "101111";
					when "011111110011100" => rgb <= "101111";
					when "011111110011101" => rgb <= "101111";
					when "011111110011110" => rgb <= "101111";
					when "011111110011111" => rgb <= "101111";
					when "100000000000000" => rgb <= "001000";
					when "100000000000001" => rgb <= "001000";
					when "100000000000010" => rgb <= "001000";
					when "100000000000011" => rgb <= "001000";
					when "100000000000100" => rgb <= "001000";
					when "100000000000101" => rgb <= "001000";
					when "100000000000110" => rgb <= "001000";
					when "100000000000111" => rgb <= "001000";
					when "100000000001000" => rgb <= "000000";
					when "100000000001001" => rgb <= "000000";
					when "100000000001010" => rgb <= "101111";
					when "100000000001011" => rgb <= "101111";
					when "100000000001100" => rgb <= "000000";
					when "100000000001101" => rgb <= "000000";
					when "100000000001110" => rgb <= "000000";
					when "100000000001111" => rgb <= "000000";
					when "100000000010000" => rgb <= "000000";
					when "100000000010001" => rgb <= "000000";
					when "100000000010010" => rgb <= "000000";
					when "100000000010011" => rgb <= "000000";
					when "100000000010100" => rgb <= "000000";
					when "100000000010101" => rgb <= "000000";
					when "100000000010110" => rgb <= "101111";
					when "100000000010111" => rgb <= "101111";
					when "100000000011000" => rgb <= "101111";
					when "100000000011001" => rgb <= "101111";
					when "100000000011010" => rgb <= "101111";
					when "100000000011011" => rgb <= "101111";
					when "100000000011100" => rgb <= "101111";
					when "100000000011101" => rgb <= "101111";
					when "100000000011110" => rgb <= "101111";
					when "100000000011111" => rgb <= "101111";
					when "100000000100000" => rgb <= "000000";
					when "100000000100001" => rgb <= "000000";
					when "100000000100010" => rgb <= "100100";
					when "100000000100011" => rgb <= "100100";
					when "100000000100100" => rgb <= "010000";
					when "100000000100101" => rgb <= "010000";
					when "100000000100110" => rgb <= "010000";
					when "100000000100111" => rgb <= "010000";
					when "100000000101000" => rgb <= "010000";
					when "100000000101001" => rgb <= "010000";
					when "100000000101010" => rgb <= "010000";
					when "100000000101011" => rgb <= "010000";
					when "100000000101100" => rgb <= "010000";
					when "100000000101101" => rgb <= "010000";
					when "100000000101110" => rgb <= "100100";
					when "100000000101111" => rgb <= "100100";
					when "100000000110000" => rgb <= "010000";
					when "100000000110001" => rgb <= "010000";
					when "100000000110010" => rgb <= "010000";
					when "100000000110011" => rgb <= "010000";
					when "100000000110100" => rgb <= "000000";
					when "100000000110101" => rgb <= "000000";
					when "100000000110110" => rgb <= "101111";
					when "100000000110111" => rgb <= "101111";
					when "100000000111000" => rgb <= "101111";
					when "100000000111001" => rgb <= "101111";
					when "100000000111010" => rgb <= "101111";
					when "100000000111011" => rgb <= "101111";
					when "100000000111100" => rgb <= "000000";
					when "100000000111101" => rgb <= "000000";
					when "100000000111110" => rgb <= "000000";
					when "100000000111111" => rgb <= "000000";
					when "100000001000000" => rgb <= "000000";
					when "100000001000001" => rgb <= "000000";
					when "100000001000010" => rgb <= "001000";
					when "100000001000011" => rgb <= "001000";
					when "100000001000100" => rgb <= "001000";
					when "100000001000101" => rgb <= "001000";
					when "100000001000110" => rgb <= "001000";
					when "100000001000111" => rgb <= "001000";
					when "100000001001000" => rgb <= "001000";
					when "100000001001001" => rgb <= "001000";
					when "100000001001010" => rgb <= "000000";
					when "100000001001011" => rgb <= "000000";
					when "100000001001100" => rgb <= "000000";
					when "100000001001101" => rgb <= "000000";
					when "100000001001110" => rgb <= "000000";
					when "100000001001111" => rgb <= "000000";
					when "100000001010000" => rgb <= "101111";
					when "100000001010001" => rgb <= "101111";
					when "100000001010010" => rgb <= "101111";
					when "100000001010011" => rgb <= "101111";
					when "100000001010100" => rgb <= "101111";
					when "100000001010101" => rgb <= "101111";
					when "100000001010110" => rgb <= "101111";
					when "100000001010111" => rgb <= "101111";
					when "100000001011000" => rgb <= "101111";
					when "100000001011001" => rgb <= "101111";
					when "100000001011010" => rgb <= "101111";
					when "100000001011011" => rgb <= "101111";
					when "100000001011100" => rgb <= "101111";
					when "100000001011101" => rgb <= "101111";
					when "100000001011110" => rgb <= "101111";
					when "100000001011111" => rgb <= "101111";
					when "100000001100000" => rgb <= "101111";
					when "100000001100001" => rgb <= "101111";
					when "100000001100010" => rgb <= "101111";
					when "100000001100011" => rgb <= "101111";
					when "100000001100100" => rgb <= "101111";
					when "100000001100101" => rgb <= "101111";
					when "100000001100110" => rgb <= "101111";
					when "100000001100111" => rgb <= "101111";
					when "100000001101000" => rgb <= "101111";
					when "100000001101001" => rgb <= "101111";
					when "100000001101010" => rgb <= "101111";
					when "100000001101011" => rgb <= "101111";
					when "100000001101100" => rgb <= "101111";
					when "100000001101101" => rgb <= "101111";
					when "100000001101110" => rgb <= "101111";
					when "100000001101111" => rgb <= "101111";
					when "100000001110000" => rgb <= "101111";
					when "100000001110001" => rgb <= "101111";
					when "100000001110010" => rgb <= "101111";
					when "100000001110011" => rgb <= "101111";
					when "100000001110100" => rgb <= "101111";
					when "100000001110101" => rgb <= "101111";
					when "100000001110110" => rgb <= "101111";
					when "100000001110111" => rgb <= "101111";
					when "100000001111000" => rgb <= "101111";
					when "100000001111001" => rgb <= "101111";
					when "100000001111010" => rgb <= "101111";
					when "100000001111011" => rgb <= "101111";
					when "100000001111100" => rgb <= "101111";
					when "100000001111101" => rgb <= "101111";
					when "100000001111110" => rgb <= "101111";
					when "100000001111111" => rgb <= "101111";
					when "100000010000000" => rgb <= "101111";
					when "100000010000001" => rgb <= "101111";
					when "100000010000010" => rgb <= "101111";
					when "100000010000011" => rgb <= "101111";
					when "100000010000100" => rgb <= "101111";
					when "100000010000101" => rgb <= "101111";
					when "100000010000110" => rgb <= "101111";
					when "100000010000111" => rgb <= "101111";
					when "100000010001000" => rgb <= "101111";
					when "100000010001001" => rgb <= "101111";
					when "100000010001010" => rgb <= "101111";
					when "100000010001011" => rgb <= "101111";
					when "100000010001100" => rgb <= "101111";
					when "100000010001101" => rgb <= "101111";
					when "100000010001110" => rgb <= "101111";
					when "100000010001111" => rgb <= "101111";
					when "100000010010000" => rgb <= "101111";
					when "100000010010001" => rgb <= "101111";
					when "100000010010010" => rgb <= "101111";
					when "100000010010011" => rgb <= "101111";
					when "100000010010100" => rgb <= "101111";
					when "100000010010101" => rgb <= "101111";
					when "100000010010110" => rgb <= "101111";
					when "100000010010111" => rgb <= "101111";
					when "100000010011000" => rgb <= "101111";
					when "100000010011001" => rgb <= "101111";
					when "100000010011010" => rgb <= "101111";
					when "100000010011011" => rgb <= "101111";
					when "100000010011100" => rgb <= "101111";
					when "100000010011101" => rgb <= "101111";
					when "100000010011110" => rgb <= "101111";
					when "100000010011111" => rgb <= "101111";
					when "100000100000000" => rgb <= "001000";
					when "100000100000001" => rgb <= "001000";
					when "100000100000010" => rgb <= "001000";
					when "100000100000011" => rgb <= "001000";
					when "100000100000100" => rgb <= "001000";
					when "100000100000101" => rgb <= "001000";
					when "100000100000110" => rgb <= "001000";
					when "100000100000111" => rgb <= "001000";
					when "100000100001000" => rgb <= "000000";
					when "100000100001001" => rgb <= "000000";
					when "100000100001010" => rgb <= "101111";
					when "100000100001011" => rgb <= "101111";
					when "100000100001100" => rgb <= "000000";
					when "100000100001101" => rgb <= "000000";
					when "100000100001110" => rgb <= "000000";
					when "100000100001111" => rgb <= "000000";
					when "100000100010000" => rgb <= "000000";
					when "100000100010001" => rgb <= "000000";
					when "100000100010010" => rgb <= "000000";
					when "100000100010011" => rgb <= "000000";
					when "100000100010100" => rgb <= "000000";
					when "100000100010101" => rgb <= "000000";
					when "100000100010110" => rgb <= "101111";
					when "100000100010111" => rgb <= "101111";
					when "100000100011000" => rgb <= "101111";
					when "100000100011001" => rgb <= "101111";
					when "100000100011010" => rgb <= "101111";
					when "100000100011011" => rgb <= "101111";
					when "100000100011100" => rgb <= "101111";
					when "100000100011101" => rgb <= "101111";
					when "100000100011110" => rgb <= "101111";
					when "100000100011111" => rgb <= "101111";
					when "100000100100000" => rgb <= "000000";
					when "100000100100001" => rgb <= "000000";
					when "100000100100010" => rgb <= "100100";
					when "100000100100011" => rgb <= "100100";
					when "100000100100100" => rgb <= "010000";
					when "100000100100101" => rgb <= "010000";
					when "100000100100110" => rgb <= "010000";
					when "100000100100111" => rgb <= "010000";
					when "100000100101000" => rgb <= "010000";
					when "100000100101001" => rgb <= "010000";
					when "100000100101010" => rgb <= "010000";
					when "100000100101011" => rgb <= "010000";
					when "100000100101100" => rgb <= "010000";
					when "100000100101101" => rgb <= "010000";
					when "100000100101110" => rgb <= "100100";
					when "100000100101111" => rgb <= "100100";
					when "100000100110000" => rgb <= "010000";
					when "100000100110001" => rgb <= "010000";
					when "100000100110010" => rgb <= "010000";
					when "100000100110011" => rgb <= "010000";
					when "100000100110100" => rgb <= "000000";
					when "100000100110101" => rgb <= "000000";
					when "100000100110110" => rgb <= "101111";
					when "100000100110111" => rgb <= "101111";
					when "100000100111000" => rgb <= "101111";
					when "100000100111001" => rgb <= "101111";
					when "100000100111010" => rgb <= "101111";
					when "100000100111011" => rgb <= "101111";
					when "100000100111100" => rgb <= "000000";
					when "100000100111101" => rgb <= "000000";
					when "100000100111110" => rgb <= "000000";
					when "100000100111111" => rgb <= "000000";
					when "100000101000000" => rgb <= "000000";
					when "100000101000001" => rgb <= "000000";
					when "100000101000010" => rgb <= "001000";
					when "100000101000011" => rgb <= "001000";
					when "100000101000100" => rgb <= "001000";
					when "100000101000101" => rgb <= "001000";
					when "100000101000110" => rgb <= "001000";
					when "100000101000111" => rgb <= "001000";
					when "100000101001000" => rgb <= "001000";
					when "100000101001001" => rgb <= "001000";
					when "100000101001010" => rgb <= "000000";
					when "100000101001011" => rgb <= "000000";
					when "100000101001100" => rgb <= "000000";
					when "100000101001101" => rgb <= "000000";
					when "100000101001110" => rgb <= "000000";
					when "100000101001111" => rgb <= "000000";
					when "100000101010000" => rgb <= "101111";
					when "100000101010001" => rgb <= "101111";
					when "100000101010010" => rgb <= "101111";
					when "100000101010011" => rgb <= "101111";
					when "100000101010100" => rgb <= "101111";
					when "100000101010101" => rgb <= "101111";
					when "100000101010110" => rgb <= "101111";
					when "100000101010111" => rgb <= "101111";
					when "100000101011000" => rgb <= "101111";
					when "100000101011001" => rgb <= "101111";
					when "100000101011010" => rgb <= "101111";
					when "100000101011011" => rgb <= "101111";
					when "100000101011100" => rgb <= "101111";
					when "100000101011101" => rgb <= "101111";
					when "100000101011110" => rgb <= "101111";
					when "100000101011111" => rgb <= "101111";
					when "100000101100000" => rgb <= "101111";
					when "100000101100001" => rgb <= "101111";
					when "100000101100010" => rgb <= "101111";
					when "100000101100011" => rgb <= "101111";
					when "100000101100100" => rgb <= "101111";
					when "100000101100101" => rgb <= "101111";
					when "100000101100110" => rgb <= "101111";
					when "100000101100111" => rgb <= "101111";
					when "100000101101000" => rgb <= "101111";
					when "100000101101001" => rgb <= "101111";
					when "100000101101010" => rgb <= "101111";
					when "100000101101011" => rgb <= "101111";
					when "100000101101100" => rgb <= "101111";
					when "100000101101101" => rgb <= "101111";
					when "100000101101110" => rgb <= "101111";
					when "100000101101111" => rgb <= "101111";
					when "100000101110000" => rgb <= "101111";
					when "100000101110001" => rgb <= "101111";
					when "100000101110010" => rgb <= "101111";
					when "100000101110011" => rgb <= "101111";
					when "100000101110100" => rgb <= "101111";
					when "100000101110101" => rgb <= "101111";
					when "100000101110110" => rgb <= "101111";
					when "100000101110111" => rgb <= "101111";
					when "100000101111000" => rgb <= "101111";
					when "100000101111001" => rgb <= "101111";
					when "100000101111010" => rgb <= "101111";
					when "100000101111011" => rgb <= "101111";
					when "100000101111100" => rgb <= "101111";
					when "100000101111101" => rgb <= "101111";
					when "100000101111110" => rgb <= "101111";
					when "100000101111111" => rgb <= "101111";
					when "100000110000000" => rgb <= "101111";
					when "100000110000001" => rgb <= "101111";
					when "100000110000010" => rgb <= "101111";
					when "100000110000011" => rgb <= "101111";
					when "100000110000100" => rgb <= "101111";
					when "100000110000101" => rgb <= "101111";
					when "100000110000110" => rgb <= "101111";
					when "100000110000111" => rgb <= "101111";
					when "100000110001000" => rgb <= "101111";
					when "100000110001001" => rgb <= "101111";
					when "100000110001010" => rgb <= "101111";
					when "100000110001011" => rgb <= "101111";
					when "100000110001100" => rgb <= "101111";
					when "100000110001101" => rgb <= "101111";
					when "100000110001110" => rgb <= "101111";
					when "100000110001111" => rgb <= "101111";
					when "100000110010000" => rgb <= "101111";
					when "100000110010001" => rgb <= "101111";
					when "100000110010010" => rgb <= "101111";
					when "100000110010011" => rgb <= "101111";
					when "100000110010100" => rgb <= "101111";
					when "100000110010101" => rgb <= "101111";
					when "100000110010110" => rgb <= "101111";
					when "100000110010111" => rgb <= "101111";
					when "100000110011000" => rgb <= "101111";
					when "100000110011001" => rgb <= "101111";
					when "100000110011010" => rgb <= "101111";
					when "100000110011011" => rgb <= "101111";
					when "100000110011100" => rgb <= "101111";
					when "100000110011101" => rgb <= "101111";
					when "100000110011110" => rgb <= "101111";
					when "100000110011111" => rgb <= "101111";
					when "100001000000000" => rgb <= "001000";
					when "100001000000001" => rgb <= "001000";
					when "100001000000010" => rgb <= "000000";
					when "100001000000011" => rgb <= "000000";
					when "100001000000100" => rgb <= "000000";
					when "100001000000101" => rgb <= "000000";
					when "100001000000110" => rgb <= "000000";
					when "100001000000111" => rgb <= "000000";
					when "100001000001000" => rgb <= "101111";
					when "100001000001001" => rgb <= "101111";
					when "100001000001010" => rgb <= "101111";
					when "100001000001011" => rgb <= "101111";
					when "100001000001100" => rgb <= "101111";
					when "100001000001101" => rgb <= "101111";
					when "100001000001110" => rgb <= "101111";
					when "100001000001111" => rgb <= "101111";
					when "100001000010000" => rgb <= "101111";
					when "100001000010001" => rgb <= "101111";
					when "100001000010010" => rgb <= "101111";
					when "100001000010011" => rgb <= "101111";
					when "100001000010100" => rgb <= "101111";
					when "100001000010101" => rgb <= "101111";
					when "100001000010110" => rgb <= "101111";
					when "100001000010111" => rgb <= "101111";
					when "100001000011000" => rgb <= "101111";
					when "100001000011001" => rgb <= "101111";
					when "100001000011010" => rgb <= "101111";
					when "100001000011011" => rgb <= "101111";
					when "100001000011100" => rgb <= "101111";
					when "100001000011101" => rgb <= "101111";
					when "100001000011110" => rgb <= "101111";
					when "100001000011111" => rgb <= "101111";
					when "100001000100000" => rgb <= "000000";
					when "100001000100001" => rgb <= "000000";
					when "100001000100010" => rgb <= "100100";
					when "100001000100011" => rgb <= "100100";
					when "100001000100100" => rgb <= "100100";
					when "100001000100101" => rgb <= "100100";
					when "100001000100110" => rgb <= "100100";
					when "100001000100111" => rgb <= "100100";
					when "100001000101000" => rgb <= "100100";
					when "100001000101001" => rgb <= "100100";
					when "100001000101010" => rgb <= "100100";
					when "100001000101011" => rgb <= "100100";
					when "100001000101100" => rgb <= "100100";
					when "100001000101101" => rgb <= "100100";
					when "100001000101110" => rgb <= "100100";
					when "100001000101111" => rgb <= "100100";
					when "100001000110000" => rgb <= "100100";
					when "100001000110001" => rgb <= "100100";
					when "100001000110010" => rgb <= "010000";
					when "100001000110011" => rgb <= "010000";
					when "100001000110100" => rgb <= "000000";
					when "100001000110101" => rgb <= "000000";
					when "100001000110110" => rgb <= "101111";
					when "100001000110111" => rgb <= "101111";
					when "100001000111000" => rgb <= "101111";
					when "100001000111001" => rgb <= "101111";
					when "100001000111010" => rgb <= "101111";
					when "100001000111011" => rgb <= "101111";
					when "100001000111100" => rgb <= "101111";
					when "100001000111101" => rgb <= "101111";
					when "100001000111110" => rgb <= "101111";
					when "100001000111111" => rgb <= "101111";
					when "100001001000000" => rgb <= "101111";
					when "100001001000001" => rgb <= "101111";
					when "100001001000010" => rgb <= "000000";
					when "100001001000011" => rgb <= "000000";
					when "100001001000100" => rgb <= "000000";
					when "100001001000101" => rgb <= "000000";
					when "100001001000110" => rgb <= "000000";
					when "100001001000111" => rgb <= "000000";
					when "100001001001000" => rgb <= "000000";
					when "100001001001001" => rgb <= "000000";
					when "100001001001010" => rgb <= "000000";
					when "100001001001011" => rgb <= "000000";
					when "100001001001100" => rgb <= "101111";
					when "100001001001101" => rgb <= "101111";
					when "100001001001110" => rgb <= "101111";
					when "100001001001111" => rgb <= "101111";
					when "100001001010000" => rgb <= "101111";
					when "100001001010001" => rgb <= "101111";
					when "100001001010010" => rgb <= "101111";
					when "100001001010011" => rgb <= "101111";
					when "100001001010100" => rgb <= "101111";
					when "100001001010101" => rgb <= "101111";
					when "100001001010110" => rgb <= "101111";
					when "100001001010111" => rgb <= "101111";
					when "100001001011000" => rgb <= "101111";
					when "100001001011001" => rgb <= "101111";
					when "100001001011010" => rgb <= "101111";
					when "100001001011011" => rgb <= "101111";
					when "100001001011100" => rgb <= "101111";
					when "100001001011101" => rgb <= "101111";
					when "100001001011110" => rgb <= "101111";
					when "100001001011111" => rgb <= "101111";
					when "100001001100000" => rgb <= "101111";
					when "100001001100001" => rgb <= "101111";
					when "100001001100010" => rgb <= "101111";
					when "100001001100011" => rgb <= "101111";
					when "100001001100100" => rgb <= "101111";
					when "100001001100101" => rgb <= "101111";
					when "100001001100110" => rgb <= "101111";
					when "100001001100111" => rgb <= "101111";
					when "100001001101000" => rgb <= "101111";
					when "100001001101001" => rgb <= "101111";
					when "100001001101010" => rgb <= "101111";
					when "100001001101011" => rgb <= "101111";
					when "100001001101100" => rgb <= "101111";
					when "100001001101101" => rgb <= "101111";
					when "100001001101110" => rgb <= "101111";
					when "100001001101111" => rgb <= "101111";
					when "100001001110000" => rgb <= "101111";
					when "100001001110001" => rgb <= "101111";
					when "100001001110010" => rgb <= "101111";
					when "100001001110011" => rgb <= "101111";
					when "100001001110100" => rgb <= "101111";
					when "100001001110101" => rgb <= "101111";
					when "100001001110110" => rgb <= "101111";
					when "100001001110111" => rgb <= "101111";
					when "100001001111000" => rgb <= "101111";
					when "100001001111001" => rgb <= "101111";
					when "100001001111010" => rgb <= "101111";
					when "100001001111011" => rgb <= "101111";
					when "100001001111100" => rgb <= "101111";
					when "100001001111101" => rgb <= "101111";
					when "100001001111110" => rgb <= "101111";
					when "100001001111111" => rgb <= "101111";
					when "100001010000000" => rgb <= "101111";
					when "100001010000001" => rgb <= "101111";
					when "100001010000010" => rgb <= "101111";
					when "100001010000011" => rgb <= "101111";
					when "100001010000100" => rgb <= "101111";
					when "100001010000101" => rgb <= "101111";
					when "100001010000110" => rgb <= "101111";
					when "100001010000111" => rgb <= "101111";
					when "100001010001000" => rgb <= "101111";
					when "100001010001001" => rgb <= "101111";
					when "100001010001010" => rgb <= "101111";
					when "100001010001011" => rgb <= "101111";
					when "100001010001100" => rgb <= "101111";
					when "100001010001101" => rgb <= "101111";
					when "100001010001110" => rgb <= "101111";
					when "100001010001111" => rgb <= "101111";
					when "100001010010000" => rgb <= "101111";
					when "100001010010001" => rgb <= "101111";
					when "100001010010010" => rgb <= "101111";
					when "100001010010011" => rgb <= "101111";
					when "100001010010100" => rgb <= "101111";
					when "100001010010101" => rgb <= "101111";
					when "100001010010110" => rgb <= "101111";
					when "100001010010111" => rgb <= "101111";
					when "100001010011000" => rgb <= "101111";
					when "100001010011001" => rgb <= "101111";
					when "100001010011010" => rgb <= "101111";
					when "100001010011011" => rgb <= "101111";
					when "100001010011100" => rgb <= "101111";
					when "100001010011101" => rgb <= "101111";
					when "100001010011110" => rgb <= "101111";
					when "100001010011111" => rgb <= "101111";
					when "100001100000000" => rgb <= "001000";
					when "100001100000001" => rgb <= "001000";
					when "100001100000010" => rgb <= "000000";
					when "100001100000011" => rgb <= "000000";
					when "100001100000100" => rgb <= "000000";
					when "100001100000101" => rgb <= "000000";
					when "100001100000110" => rgb <= "000000";
					when "100001100000111" => rgb <= "000000";
					when "100001100001000" => rgb <= "101111";
					when "100001100001001" => rgb <= "101111";
					when "100001100001010" => rgb <= "101111";
					when "100001100001011" => rgb <= "101111";
					when "100001100001100" => rgb <= "101111";
					when "100001100001101" => rgb <= "101111";
					when "100001100001110" => rgb <= "101111";
					when "100001100001111" => rgb <= "101111";
					when "100001100010000" => rgb <= "101111";
					when "100001100010001" => rgb <= "101111";
					when "100001100010010" => rgb <= "101111";
					when "100001100010011" => rgb <= "101111";
					when "100001100010100" => rgb <= "101111";
					when "100001100010101" => rgb <= "101111";
					when "100001100010110" => rgb <= "101111";
					when "100001100010111" => rgb <= "101111";
					when "100001100011000" => rgb <= "101111";
					when "100001100011001" => rgb <= "101111";
					when "100001100011010" => rgb <= "101111";
					when "100001100011011" => rgb <= "101111";
					when "100001100011100" => rgb <= "101111";
					when "100001100011101" => rgb <= "101111";
					when "100001100011110" => rgb <= "101111";
					when "100001100011111" => rgb <= "101111";
					when "100001100100000" => rgb <= "000000";
					when "100001100100001" => rgb <= "000000";
					when "100001100100010" => rgb <= "100100";
					when "100001100100011" => rgb <= "100100";
					when "100001100100100" => rgb <= "100100";
					when "100001100100101" => rgb <= "100100";
					when "100001100100110" => rgb <= "100100";
					when "100001100100111" => rgb <= "100100";
					when "100001100101000" => rgb <= "100100";
					when "100001100101001" => rgb <= "100100";
					when "100001100101010" => rgb <= "100100";
					when "100001100101011" => rgb <= "100100";
					when "100001100101100" => rgb <= "100100";
					when "100001100101101" => rgb <= "100100";
					when "100001100101110" => rgb <= "100100";
					when "100001100101111" => rgb <= "100100";
					when "100001100110000" => rgb <= "100100";
					when "100001100110001" => rgb <= "100100";
					when "100001100110010" => rgb <= "010000";
					when "100001100110011" => rgb <= "010000";
					when "100001100110100" => rgb <= "000000";
					when "100001100110101" => rgb <= "000000";
					when "100001100110110" => rgb <= "101111";
					when "100001100110111" => rgb <= "101111";
					when "100001100111000" => rgb <= "101111";
					when "100001100111001" => rgb <= "101111";
					when "100001100111010" => rgb <= "101111";
					when "100001100111011" => rgb <= "101111";
					when "100001100111100" => rgb <= "101111";
					when "100001100111101" => rgb <= "101111";
					when "100001100111110" => rgb <= "101111";
					when "100001100111111" => rgb <= "101111";
					when "100001101000000" => rgb <= "101111";
					when "100001101000001" => rgb <= "101111";
					when "100001101000010" => rgb <= "000000";
					when "100001101000011" => rgb <= "000000";
					when "100001101000100" => rgb <= "000000";
					when "100001101000101" => rgb <= "000000";
					when "100001101000110" => rgb <= "000000";
					when "100001101000111" => rgb <= "000000";
					when "100001101001000" => rgb <= "000000";
					when "100001101001001" => rgb <= "000000";
					when "100001101001010" => rgb <= "000000";
					when "100001101001011" => rgb <= "000000";
					when "100001101001100" => rgb <= "101111";
					when "100001101001101" => rgb <= "101111";
					when "100001101001110" => rgb <= "101111";
					when "100001101001111" => rgb <= "101111";
					when "100001101010000" => rgb <= "101111";
					when "100001101010001" => rgb <= "101111";
					when "100001101010010" => rgb <= "101111";
					when "100001101010011" => rgb <= "101111";
					when "100001101010100" => rgb <= "101111";
					when "100001101010101" => rgb <= "101111";
					when "100001101010110" => rgb <= "101111";
					when "100001101010111" => rgb <= "101111";
					when "100001101011000" => rgb <= "101111";
					when "100001101011001" => rgb <= "101111";
					when "100001101011010" => rgb <= "101111";
					when "100001101011011" => rgb <= "101111";
					when "100001101011100" => rgb <= "101111";
					when "100001101011101" => rgb <= "101111";
					when "100001101011110" => rgb <= "101111";
					when "100001101011111" => rgb <= "101111";
					when "100001101100000" => rgb <= "101111";
					when "100001101100001" => rgb <= "101111";
					when "100001101100010" => rgb <= "101111";
					when "100001101100011" => rgb <= "101111";
					when "100001101100100" => rgb <= "101111";
					when "100001101100101" => rgb <= "101111";
					when "100001101100110" => rgb <= "101111";
					when "100001101100111" => rgb <= "101111";
					when "100001101101000" => rgb <= "101111";
					when "100001101101001" => rgb <= "101111";
					when "100001101101010" => rgb <= "101111";
					when "100001101101011" => rgb <= "101111";
					when "100001101101100" => rgb <= "101111";
					when "100001101101101" => rgb <= "101111";
					when "100001101101110" => rgb <= "101111";
					when "100001101101111" => rgb <= "101111";
					when "100001101110000" => rgb <= "101111";
					when "100001101110001" => rgb <= "101111";
					when "100001101110010" => rgb <= "101111";
					when "100001101110011" => rgb <= "101111";
					when "100001101110100" => rgb <= "101111";
					when "100001101110101" => rgb <= "101111";
					when "100001101110110" => rgb <= "101111";
					when "100001101110111" => rgb <= "101111";
					when "100001101111000" => rgb <= "101111";
					when "100001101111001" => rgb <= "101111";
					when "100001101111010" => rgb <= "101111";
					when "100001101111011" => rgb <= "101111";
					when "100001101111100" => rgb <= "101111";
					when "100001101111101" => rgb <= "101111";
					when "100001101111110" => rgb <= "101111";
					when "100001101111111" => rgb <= "101111";
					when "100001110000000" => rgb <= "101111";
					when "100001110000001" => rgb <= "101111";
					when "100001110000010" => rgb <= "101111";
					when "100001110000011" => rgb <= "101111";
					when "100001110000100" => rgb <= "101111";
					when "100001110000101" => rgb <= "101111";
					when "100001110000110" => rgb <= "101111";
					when "100001110000111" => rgb <= "101111";
					when "100001110001000" => rgb <= "101111";
					when "100001110001001" => rgb <= "101111";
					when "100001110001010" => rgb <= "101111";
					when "100001110001011" => rgb <= "101111";
					when "100001110001100" => rgb <= "101111";
					when "100001110001101" => rgb <= "101111";
					when "100001110001110" => rgb <= "101111";
					when "100001110001111" => rgb <= "101111";
					when "100001110010000" => rgb <= "101111";
					when "100001110010001" => rgb <= "101111";
					when "100001110010010" => rgb <= "101111";
					when "100001110010011" => rgb <= "101111";
					when "100001110010100" => rgb <= "101111";
					when "100001110010101" => rgb <= "101111";
					when "100001110010110" => rgb <= "101111";
					when "100001110010111" => rgb <= "101111";
					when "100001110011000" => rgb <= "101111";
					when "100001110011001" => rgb <= "101111";
					when "100001110011010" => rgb <= "101111";
					when "100001110011011" => rgb <= "101111";
					when "100001110011100" => rgb <= "101111";
					when "100001110011101" => rgb <= "101111";
					when "100001110011110" => rgb <= "101111";
					when "100001110011111" => rgb <= "101111";
					when "100010000000000" => rgb <= "000000";
					when "100010000000001" => rgb <= "000000";
					when "100010000000010" => rgb <= "000000";
					when "100010000000011" => rgb <= "000000";
					when "100010000000100" => rgb <= "101111";
					when "100010000000101" => rgb <= "101111";
					when "100010000000110" => rgb <= "101111";
					when "100010000000111" => rgb <= "101111";
					when "100010000001000" => rgb <= "101111";
					when "100010000001001" => rgb <= "101111";
					when "100010000001010" => rgb <= "101111";
					when "100010000001011" => rgb <= "101111";
					when "100010000001100" => rgb <= "101111";
					when "100010000001101" => rgb <= "101111";
					when "100010000001110" => rgb <= "101111";
					when "100010000001111" => rgb <= "101111";
					when "100010000010000" => rgb <= "101111";
					when "100010000010001" => rgb <= "101111";
					when "100010000010010" => rgb <= "101111";
					when "100010000010011" => rgb <= "101111";
					when "100010000010100" => rgb <= "101111";
					when "100010000010101" => rgb <= "101111";
					when "100010000010110" => rgb <= "101111";
					when "100010000010111" => rgb <= "101111";
					when "100010000011000" => rgb <= "101111";
					when "100010000011001" => rgb <= "101111";
					when "100010000011010" => rgb <= "101111";
					when "100010000011011" => rgb <= "101111";
					when "100010000011100" => rgb <= "101111";
					when "100010000011101" => rgb <= "101111";
					when "100010000011110" => rgb <= "101111";
					when "100010000011111" => rgb <= "101111";
					when "100010000100000" => rgb <= "000000";
					when "100010000100001" => rgb <= "000000";
					when "100010000100010" => rgb <= "100100";
					when "100010000100011" => rgb <= "100100";
					when "100010000100100" => rgb <= "100100";
					when "100010000100101" => rgb <= "100100";
					when "100010000100110" => rgb <= "100100";
					when "100010000100111" => rgb <= "100100";
					when "100010000101000" => rgb <= "000000";
					when "100010000101001" => rgb <= "000000";
					when "100010000101010" => rgb <= "100100";
					when "100010000101011" => rgb <= "100100";
					when "100010000101100" => rgb <= "100100";
					when "100010000101101" => rgb <= "100100";
					when "100010000101110" => rgb <= "100100";
					when "100010000101111" => rgb <= "100100";
					when "100010000110000" => rgb <= "000000";
					when "100010000110001" => rgb <= "000000";
					when "100010000110010" => rgb <= "010000";
					when "100010000110011" => rgb <= "010000";
					when "100010000110100" => rgb <= "000000";
					when "100010000110101" => rgb <= "000000";
					when "100010000110110" => rgb <= "101111";
					when "100010000110111" => rgb <= "101111";
					when "100010000111000" => rgb <= "101111";
					when "100010000111001" => rgb <= "101111";
					when "100010000111010" => rgb <= "101111";
					when "100010000111011" => rgb <= "101111";
					when "100010000111100" => rgb <= "101111";
					when "100010000111101" => rgb <= "101111";
					when "100010000111110" => rgb <= "101111";
					when "100010000111111" => rgb <= "101111";
					when "100010001000000" => rgb <= "101111";
					when "100010001000001" => rgb <= "101111";
					when "100010001000010" => rgb <= "101111";
					when "100010001000011" => rgb <= "101111";
					when "100010001000100" => rgb <= "101111";
					when "100010001000101" => rgb <= "101111";
					when "100010001000110" => rgb <= "000000";
					when "100010001000111" => rgb <= "000000";
					when "100010001001000" => rgb <= "101111";
					when "100010001001001" => rgb <= "101111";
					when "100010001001010" => rgb <= "101111";
					when "100010001001011" => rgb <= "101111";
					when "100010001001100" => rgb <= "101111";
					when "100010001001101" => rgb <= "101111";
					when "100010001001110" => rgb <= "101111";
					when "100010001001111" => rgb <= "101111";
					when "100010001010000" => rgb <= "101111";
					when "100010001010001" => rgb <= "101111";
					when "100010001010010" => rgb <= "101111";
					when "100010001010011" => rgb <= "101111";
					when "100010001010100" => rgb <= "101111";
					when "100010001010101" => rgb <= "101111";
					when "100010001010110" => rgb <= "101111";
					when "100010001010111" => rgb <= "101111";
					when "100010001011000" => rgb <= "101111";
					when "100010001011001" => rgb <= "101111";
					when "100010001011010" => rgb <= "101111";
					when "100010001011011" => rgb <= "101111";
					when "100010001011100" => rgb <= "101111";
					when "100010001011101" => rgb <= "101111";
					when "100010001011110" => rgb <= "101111";
					when "100010001011111" => rgb <= "101111";
					when "100010001100000" => rgb <= "101111";
					when "100010001100001" => rgb <= "101111";
					when "100010001100010" => rgb <= "101111";
					when "100010001100011" => rgb <= "101111";
					when "100010001100100" => rgb <= "101111";
					when "100010001100101" => rgb <= "101111";
					when "100010001100110" => rgb <= "101111";
					when "100010001100111" => rgb <= "101111";
					when "100010001101000" => rgb <= "101111";
					when "100010001101001" => rgb <= "101111";
					when "100010001101010" => rgb <= "101111";
					when "100010001101011" => rgb <= "101111";
					when "100010001101100" => rgb <= "101111";
					when "100010001101101" => rgb <= "101111";
					when "100010001101110" => rgb <= "101111";
					when "100010001101111" => rgb <= "101111";
					when "100010001110000" => rgb <= "101111";
					when "100010001110001" => rgb <= "101111";
					when "100010001110010" => rgb <= "101111";
					when "100010001110011" => rgb <= "101111";
					when "100010001110100" => rgb <= "101111";
					when "100010001110101" => rgb <= "101111";
					when "100010001110110" => rgb <= "101111";
					when "100010001110111" => rgb <= "101111";
					when "100010001111000" => rgb <= "101111";
					when "100010001111001" => rgb <= "101111";
					when "100010001111010" => rgb <= "101111";
					when "100010001111011" => rgb <= "101111";
					when "100010001111100" => rgb <= "101111";
					when "100010001111101" => rgb <= "101111";
					when "100010001111110" => rgb <= "101111";
					when "100010001111111" => rgb <= "101111";
					when "100010010000000" => rgb <= "101111";
					when "100010010000001" => rgb <= "101111";
					when "100010010000010" => rgb <= "101111";
					when "100010010000011" => rgb <= "101111";
					when "100010010000100" => rgb <= "101111";
					when "100010010000101" => rgb <= "101111";
					when "100010010000110" => rgb <= "101111";
					when "100010010000111" => rgb <= "101111";
					when "100010010001000" => rgb <= "101111";
					when "100010010001001" => rgb <= "101111";
					when "100010010001010" => rgb <= "101111";
					when "100010010001011" => rgb <= "101111";
					when "100010010001100" => rgb <= "101111";
					when "100010010001101" => rgb <= "101111";
					when "100010010001110" => rgb <= "101111";
					when "100010010001111" => rgb <= "101111";
					when "100010010010000" => rgb <= "101111";
					when "100010010010001" => rgb <= "101111";
					when "100010010010010" => rgb <= "101111";
					when "100010010010011" => rgb <= "101111";
					when "100010010010100" => rgb <= "101111";
					when "100010010010101" => rgb <= "101111";
					when "100010010010110" => rgb <= "101111";
					when "100010010010111" => rgb <= "101111";
					when "100010010011000" => rgb <= "101111";
					when "100010010011001" => rgb <= "101111";
					when "100010010011010" => rgb <= "101111";
					when "100010010011011" => rgb <= "101111";
					when "100010010011100" => rgb <= "101111";
					when "100010010011101" => rgb <= "101111";
					when "100010010011110" => rgb <= "101111";
					when "100010010011111" => rgb <= "101111";
					when "100010100000000" => rgb <= "000000";
					when "100010100000001" => rgb <= "000000";
					when "100010100000010" => rgb <= "000000";
					when "100010100000011" => rgb <= "000000";
					when "100010100000100" => rgb <= "101111";
					when "100010100000101" => rgb <= "101111";
					when "100010100000110" => rgb <= "101111";
					when "100010100000111" => rgb <= "101111";
					when "100010100001000" => rgb <= "101111";
					when "100010100001001" => rgb <= "101111";
					when "100010100001010" => rgb <= "101111";
					when "100010100001011" => rgb <= "101111";
					when "100010100001100" => rgb <= "101111";
					when "100010100001101" => rgb <= "101111";
					when "100010100001110" => rgb <= "101111";
					when "100010100001111" => rgb <= "101111";
					when "100010100010000" => rgb <= "101111";
					when "100010100010001" => rgb <= "101111";
					when "100010100010010" => rgb <= "101111";
					when "100010100010011" => rgb <= "101111";
					when "100010100010100" => rgb <= "101111";
					when "100010100010101" => rgb <= "101111";
					when "100010100010110" => rgb <= "101111";
					when "100010100010111" => rgb <= "101111";
					when "100010100011000" => rgb <= "101111";
					when "100010100011001" => rgb <= "101111";
					when "100010100011010" => rgb <= "101111";
					when "100010100011011" => rgb <= "101111";
					when "100010100011100" => rgb <= "101111";
					when "100010100011101" => rgb <= "101111";
					when "100010100011110" => rgb <= "101111";
					when "100010100011111" => rgb <= "101111";
					when "100010100100000" => rgb <= "000000";
					when "100010100100001" => rgb <= "000000";
					when "100010100100010" => rgb <= "100100";
					when "100010100100011" => rgb <= "100100";
					when "100010100100100" => rgb <= "100100";
					when "100010100100101" => rgb <= "100100";
					when "100010100100110" => rgb <= "100100";
					when "100010100100111" => rgb <= "100100";
					when "100010100101000" => rgb <= "000000";
					when "100010100101001" => rgb <= "000000";
					when "100010100101010" => rgb <= "100100";
					when "100010100101011" => rgb <= "100100";
					when "100010100101100" => rgb <= "100100";
					when "100010100101101" => rgb <= "100100";
					when "100010100101110" => rgb <= "100100";
					when "100010100101111" => rgb <= "100100";
					when "100010100110000" => rgb <= "000000";
					when "100010100110001" => rgb <= "000000";
					when "100010100110010" => rgb <= "010000";
					when "100010100110011" => rgb <= "010000";
					when "100010100110100" => rgb <= "000000";
					when "100010100110101" => rgb <= "000000";
					when "100010100110110" => rgb <= "101111";
					when "100010100110111" => rgb <= "101111";
					when "100010100111000" => rgb <= "101111";
					when "100010100111001" => rgb <= "101111";
					when "100010100111010" => rgb <= "101111";
					when "100010100111011" => rgb <= "101111";
					when "100010100111100" => rgb <= "101111";
					when "100010100111101" => rgb <= "101111";
					when "100010100111110" => rgb <= "101111";
					when "100010100111111" => rgb <= "101111";
					when "100010101000000" => rgb <= "101111";
					when "100010101000001" => rgb <= "101111";
					when "100010101000010" => rgb <= "101111";
					when "100010101000011" => rgb <= "101111";
					when "100010101000100" => rgb <= "101111";
					when "100010101000101" => rgb <= "101111";
					when "100010101000110" => rgb <= "000000";
					when "100010101000111" => rgb <= "000000";
					when "100010101001000" => rgb <= "101111";
					when "100010101001001" => rgb <= "101111";
					when "100010101001010" => rgb <= "101111";
					when "100010101001011" => rgb <= "101111";
					when "100010101001100" => rgb <= "101111";
					when "100010101001101" => rgb <= "101111";
					when "100010101001110" => rgb <= "101111";
					when "100010101001111" => rgb <= "101111";
					when "100010101010000" => rgb <= "101111";
					when "100010101010001" => rgb <= "101111";
					when "100010101010010" => rgb <= "101111";
					when "100010101010011" => rgb <= "101111";
					when "100010101010100" => rgb <= "101111";
					when "100010101010101" => rgb <= "101111";
					when "100010101010110" => rgb <= "101111";
					when "100010101010111" => rgb <= "101111";
					when "100010101011000" => rgb <= "101111";
					when "100010101011001" => rgb <= "101111";
					when "100010101011010" => rgb <= "101111";
					when "100010101011011" => rgb <= "101111";
					when "100010101011100" => rgb <= "101111";
					when "100010101011101" => rgb <= "101111";
					when "100010101011110" => rgb <= "101111";
					when "100010101011111" => rgb <= "101111";
					when "100010101100000" => rgb <= "101111";
					when "100010101100001" => rgb <= "101111";
					when "100010101100010" => rgb <= "101111";
					when "100010101100011" => rgb <= "101111";
					when "100010101100100" => rgb <= "101111";
					when "100010101100101" => rgb <= "101111";
					when "100010101100110" => rgb <= "101111";
					when "100010101100111" => rgb <= "101111";
					when "100010101101000" => rgb <= "101111";
					when "100010101101001" => rgb <= "101111";
					when "100010101101010" => rgb <= "101111";
					when "100010101101011" => rgb <= "101111";
					when "100010101101100" => rgb <= "101111";
					when "100010101101101" => rgb <= "101111";
					when "100010101101110" => rgb <= "101111";
					when "100010101101111" => rgb <= "101111";
					when "100010101110000" => rgb <= "101111";
					when "100010101110001" => rgb <= "101111";
					when "100010101110010" => rgb <= "101111";
					when "100010101110011" => rgb <= "101111";
					when "100010101110100" => rgb <= "101111";
					when "100010101110101" => rgb <= "101111";
					when "100010101110110" => rgb <= "101111";
					when "100010101110111" => rgb <= "101111";
					when "100010101111000" => rgb <= "101111";
					when "100010101111001" => rgb <= "101111";
					when "100010101111010" => rgb <= "101111";
					when "100010101111011" => rgb <= "101111";
					when "100010101111100" => rgb <= "101111";
					when "100010101111101" => rgb <= "101111";
					when "100010101111110" => rgb <= "101111";
					when "100010101111111" => rgb <= "101111";
					when "100010110000000" => rgb <= "101111";
					when "100010110000001" => rgb <= "101111";
					when "100010110000010" => rgb <= "101111";
					when "100010110000011" => rgb <= "101111";
					when "100010110000100" => rgb <= "101111";
					when "100010110000101" => rgb <= "101111";
					when "100010110000110" => rgb <= "101111";
					when "100010110000111" => rgb <= "101111";
					when "100010110001000" => rgb <= "101111";
					when "100010110001001" => rgb <= "101111";
					when "100010110001010" => rgb <= "101111";
					when "100010110001011" => rgb <= "101111";
					when "100010110001100" => rgb <= "101111";
					when "100010110001101" => rgb <= "101111";
					when "100010110001110" => rgb <= "101111";
					when "100010110001111" => rgb <= "101111";
					when "100010110010000" => rgb <= "101111";
					when "100010110010001" => rgb <= "101111";
					when "100010110010010" => rgb <= "101111";
					when "100010110010011" => rgb <= "101111";
					when "100010110010100" => rgb <= "101111";
					when "100010110010101" => rgb <= "101111";
					when "100010110010110" => rgb <= "101111";
					when "100010110010111" => rgb <= "101111";
					when "100010110011000" => rgb <= "101111";
					when "100010110011001" => rgb <= "101111";
					when "100010110011010" => rgb <= "101111";
					when "100010110011011" => rgb <= "101111";
					when "100010110011100" => rgb <= "101111";
					when "100010110011101" => rgb <= "101111";
					when "100010110011110" => rgb <= "101111";
					when "100010110011111" => rgb <= "101111";
					when "100011000000000" => rgb <= "101111";
					when "100011000000001" => rgb <= "101111";
					when "100011000000010" => rgb <= "101111";
					when "100011000000011" => rgb <= "101111";
					when "100011000000100" => rgb <= "101111";
					when "100011000000101" => rgb <= "101111";
					when "100011000000110" => rgb <= "101111";
					when "100011000000111" => rgb <= "101111";
					when "100011000001000" => rgb <= "101111";
					when "100011000001001" => rgb <= "101111";
					when "100011000001010" => rgb <= "101111";
					when "100011000001011" => rgb <= "101111";
					when "100011000001100" => rgb <= "101111";
					when "100011000001101" => rgb <= "101111";
					when "100011000001110" => rgb <= "101111";
					when "100011000001111" => rgb <= "101111";
					when "100011000010000" => rgb <= "101111";
					when "100011000010001" => rgb <= "101111";
					when "100011000010010" => rgb <= "101111";
					when "100011000010011" => rgb <= "101111";
					when "100011000010100" => rgb <= "101111";
					when "100011000010101" => rgb <= "101111";
					when "100011000010110" => rgb <= "101111";
					when "100011000010111" => rgb <= "101111";
					when "100011000011000" => rgb <= "101111";
					when "100011000011001" => rgb <= "101111";
					when "100011000011010" => rgb <= "101111";
					when "100011000011011" => rgb <= "101111";
					when "100011000011100" => rgb <= "101111";
					when "100011000011101" => rgb <= "101111";
					when "100011000011110" => rgb <= "101111";
					when "100011000011111" => rgb <= "101111";
					when "100011000100000" => rgb <= "000000";
					when "100011000100001" => rgb <= "000000";
					when "100011000100010" => rgb <= "100100";
					when "100011000100011" => rgb <= "100100";
					when "100011000100100" => rgb <= "100100";
					when "100011000100101" => rgb <= "100100";
					when "100011000100110" => rgb <= "000000";
					when "100011000100111" => rgb <= "000000";
					when "100011000101000" => rgb <= "000000";
					when "100011000101001" => rgb <= "000000";
					when "100011000101010" => rgb <= "000000";
					when "100011000101011" => rgb <= "000000";
					when "100011000101100" => rgb <= "100100";
					when "100011000101101" => rgb <= "100100";
					when "100011000101110" => rgb <= "000000";
					when "100011000101111" => rgb <= "000000";
					when "100011000110000" => rgb <= "000000";
					when "100011000110001" => rgb <= "000000";
					when "100011000110010" => rgb <= "000000";
					when "100011000110011" => rgb <= "000000";
					when "100011000110100" => rgb <= "000000";
					when "100011000110101" => rgb <= "000000";
					when "100011000110110" => rgb <= "101111";
					when "100011000110111" => rgb <= "101111";
					when "100011000111000" => rgb <= "101111";
					when "100011000111001" => rgb <= "101111";
					when "100011000111010" => rgb <= "101111";
					when "100011000111011" => rgb <= "101111";
					when "100011000111100" => rgb <= "101111";
					when "100011000111101" => rgb <= "101111";
					when "100011000111110" => rgb <= "101111";
					when "100011000111111" => rgb <= "101111";
					when "100011001000000" => rgb <= "101111";
					when "100011001000001" => rgb <= "101111";
					when "100011001000010" => rgb <= "101111";
					when "100011001000011" => rgb <= "101111";
					when "100011001000100" => rgb <= "101111";
					when "100011001000101" => rgb <= "101111";
					when "100011001000110" => rgb <= "101111";
					when "100011001000111" => rgb <= "101111";
					when "100011001001000" => rgb <= "101111";
					when "100011001001001" => rgb <= "101111";
					when "100011001001010" => rgb <= "101111";
					when "100011001001011" => rgb <= "101111";
					when "100011001001100" => rgb <= "101111";
					when "100011001001101" => rgb <= "101111";
					when "100011001001110" => rgb <= "101111";
					when "100011001001111" => rgb <= "101111";
					when "100011001010000" => rgb <= "101111";
					when "100011001010001" => rgb <= "101111";
					when "100011001010010" => rgb <= "101111";
					when "100011001010011" => rgb <= "101111";
					when "100011001010100" => rgb <= "101111";
					when "100011001010101" => rgb <= "101111";
					when "100011001010110" => rgb <= "101111";
					when "100011001010111" => rgb <= "101111";
					when "100011001011000" => rgb <= "101111";
					when "100011001011001" => rgb <= "101111";
					when "100011001011010" => rgb <= "101111";
					when "100011001011011" => rgb <= "101111";
					when "100011001011100" => rgb <= "101111";
					when "100011001011101" => rgb <= "101111";
					when "100011001011110" => rgb <= "101111";
					when "100011001011111" => rgb <= "101111";
					when "100011001100000" => rgb <= "101111";
					when "100011001100001" => rgb <= "101111";
					when "100011001100010" => rgb <= "101111";
					when "100011001100011" => rgb <= "101111";
					when "100011001100100" => rgb <= "101111";
					when "100011001100101" => rgb <= "101111";
					when "100011001100110" => rgb <= "101111";
					when "100011001100111" => rgb <= "101111";
					when "100011001101000" => rgb <= "101111";
					when "100011001101001" => rgb <= "101111";
					when "100011001101010" => rgb <= "101111";
					when "100011001101011" => rgb <= "101111";
					when "100011001101100" => rgb <= "101111";
					when "100011001101101" => rgb <= "101111";
					when "100011001101110" => rgb <= "101111";
					when "100011001101111" => rgb <= "101111";
					when "100011001110000" => rgb <= "101111";
					when "100011001110001" => rgb <= "101111";
					when "100011001110010" => rgb <= "101111";
					when "100011001110011" => rgb <= "101111";
					when "100011001110100" => rgb <= "101111";
					when "100011001110101" => rgb <= "101111";
					when "100011001110110" => rgb <= "101111";
					when "100011001110111" => rgb <= "101111";
					when "100011001111000" => rgb <= "101111";
					when "100011001111001" => rgb <= "101111";
					when "100011001111010" => rgb <= "101111";
					when "100011001111011" => rgb <= "101111";
					when "100011001111100" => rgb <= "101111";
					when "100011001111101" => rgb <= "101111";
					when "100011001111110" => rgb <= "101111";
					when "100011001111111" => rgb <= "101111";
					when "100011010000000" => rgb <= "101111";
					when "100011010000001" => rgb <= "101111";
					when "100011010000010" => rgb <= "101111";
					when "100011010000011" => rgb <= "101111";
					when "100011010000100" => rgb <= "101111";
					when "100011010000101" => rgb <= "101111";
					when "100011010000110" => rgb <= "101111";
					when "100011010000111" => rgb <= "101111";
					when "100011010001000" => rgb <= "101111";
					when "100011010001001" => rgb <= "101111";
					when "100011010001010" => rgb <= "101111";
					when "100011010001011" => rgb <= "101111";
					when "100011010001100" => rgb <= "101111";
					when "100011010001101" => rgb <= "101111";
					when "100011010001110" => rgb <= "101111";
					when "100011010001111" => rgb <= "101111";
					when "100011010010000" => rgb <= "101111";
					when "100011010010001" => rgb <= "101111";
					when "100011010010010" => rgb <= "101111";
					when "100011010010011" => rgb <= "101111";
					when "100011010010100" => rgb <= "101111";
					when "100011010010101" => rgb <= "101111";
					when "100011010010110" => rgb <= "101111";
					when "100011010010111" => rgb <= "101111";
					when "100011010011000" => rgb <= "101111";
					when "100011010011001" => rgb <= "101111";
					when "100011010011010" => rgb <= "101111";
					when "100011010011011" => rgb <= "101111";
					when "100011010011100" => rgb <= "101111";
					when "100011010011101" => rgb <= "101111";
					when "100011010011110" => rgb <= "101111";
					when "100011010011111" => rgb <= "101111";
					when "100011100000000" => rgb <= "101111";
					when "100011100000001" => rgb <= "101111";
					when "100011100000010" => rgb <= "101111";
					when "100011100000011" => rgb <= "101111";
					when "100011100000100" => rgb <= "101111";
					when "100011100000101" => rgb <= "101111";
					when "100011100000110" => rgb <= "101111";
					when "100011100000111" => rgb <= "101111";
					when "100011100001000" => rgb <= "101111";
					when "100011100001001" => rgb <= "101111";
					when "100011100001010" => rgb <= "101111";
					when "100011100001011" => rgb <= "101111";
					when "100011100001100" => rgb <= "101111";
					when "100011100001101" => rgb <= "101111";
					when "100011100001110" => rgb <= "101111";
					when "100011100001111" => rgb <= "101111";
					when "100011100010000" => rgb <= "101111";
					when "100011100010001" => rgb <= "101111";
					when "100011100010010" => rgb <= "101111";
					when "100011100010011" => rgb <= "101111";
					when "100011100010100" => rgb <= "101111";
					when "100011100010101" => rgb <= "101111";
					when "100011100010110" => rgb <= "101111";
					when "100011100010111" => rgb <= "101111";
					when "100011100011000" => rgb <= "101111";
					when "100011100011001" => rgb <= "101111";
					when "100011100011010" => rgb <= "101111";
					when "100011100011011" => rgb <= "101111";
					when "100011100011100" => rgb <= "101111";
					when "100011100011101" => rgb <= "101111";
					when "100011100011110" => rgb <= "101111";
					when "100011100011111" => rgb <= "101111";
					when "100011100100000" => rgb <= "000000";
					when "100011100100001" => rgb <= "000000";
					when "100011100100010" => rgb <= "100100";
					when "100011100100011" => rgb <= "100100";
					when "100011100100100" => rgb <= "100100";
					when "100011100100101" => rgb <= "100100";
					when "100011100100110" => rgb <= "000000";
					when "100011100100111" => rgb <= "000000";
					when "100011100101000" => rgb <= "000000";
					when "100011100101001" => rgb <= "000000";
					when "100011100101010" => rgb <= "000000";
					when "100011100101011" => rgb <= "000000";
					when "100011100101100" => rgb <= "100100";
					when "100011100101101" => rgb <= "100100";
					when "100011100101110" => rgb <= "000000";
					when "100011100101111" => rgb <= "000000";
					when "100011100110000" => rgb <= "000000";
					when "100011100110001" => rgb <= "000000";
					when "100011100110010" => rgb <= "000000";
					when "100011100110011" => rgb <= "000000";
					when "100011100110100" => rgb <= "000000";
					when "100011100110101" => rgb <= "000000";
					when "100011100110110" => rgb <= "101111";
					when "100011100110111" => rgb <= "101111";
					when "100011100111000" => rgb <= "101111";
					when "100011100111001" => rgb <= "101111";
					when "100011100111010" => rgb <= "101111";
					when "100011100111011" => rgb <= "101111";
					when "100011100111100" => rgb <= "101111";
					when "100011100111101" => rgb <= "101111";
					when "100011100111110" => rgb <= "101111";
					when "100011100111111" => rgb <= "101111";
					when "100011101000000" => rgb <= "101111";
					when "100011101000001" => rgb <= "101111";
					when "100011101000010" => rgb <= "101111";
					when "100011101000011" => rgb <= "101111";
					when "100011101000100" => rgb <= "101111";
					when "100011101000101" => rgb <= "101111";
					when "100011101000110" => rgb <= "101111";
					when "100011101000111" => rgb <= "101111";
					when "100011101001000" => rgb <= "101111";
					when "100011101001001" => rgb <= "101111";
					when "100011101001010" => rgb <= "101111";
					when "100011101001011" => rgb <= "101111";
					when "100011101001100" => rgb <= "101111";
					when "100011101001101" => rgb <= "101111";
					when "100011101001110" => rgb <= "101111";
					when "100011101001111" => rgb <= "101111";
					when "100011101010000" => rgb <= "101111";
					when "100011101010001" => rgb <= "101111";
					when "100011101010010" => rgb <= "101111";
					when "100011101010011" => rgb <= "101111";
					when "100011101010100" => rgb <= "101111";
					when "100011101010101" => rgb <= "101111";
					when "100011101010110" => rgb <= "101111";
					when "100011101010111" => rgb <= "101111";
					when "100011101011000" => rgb <= "101111";
					when "100011101011001" => rgb <= "101111";
					when "100011101011010" => rgb <= "101111";
					when "100011101011011" => rgb <= "101111";
					when "100011101011100" => rgb <= "101111";
					when "100011101011101" => rgb <= "101111";
					when "100011101011110" => rgb <= "101111";
					when "100011101011111" => rgb <= "101111";
					when "100011101100000" => rgb <= "101111";
					when "100011101100001" => rgb <= "101111";
					when "100011101100010" => rgb <= "101111";
					when "100011101100011" => rgb <= "101111";
					when "100011101100100" => rgb <= "101111";
					when "100011101100101" => rgb <= "101111";
					when "100011101100110" => rgb <= "101111";
					when "100011101100111" => rgb <= "101111";
					when "100011101101000" => rgb <= "101111";
					when "100011101101001" => rgb <= "101111";
					when "100011101101010" => rgb <= "101111";
					when "100011101101011" => rgb <= "101111";
					when "100011101101100" => rgb <= "101111";
					when "100011101101101" => rgb <= "101111";
					when "100011101101110" => rgb <= "101111";
					when "100011101101111" => rgb <= "101111";
					when "100011101110000" => rgb <= "101111";
					when "100011101110001" => rgb <= "101111";
					when "100011101110010" => rgb <= "101111";
					when "100011101110011" => rgb <= "101111";
					when "100011101110100" => rgb <= "101111";
					when "100011101110101" => rgb <= "101111";
					when "100011101110110" => rgb <= "101111";
					when "100011101110111" => rgb <= "101111";
					when "100011101111000" => rgb <= "101111";
					when "100011101111001" => rgb <= "101111";
					when "100011101111010" => rgb <= "101111";
					when "100011101111011" => rgb <= "101111";
					when "100011101111100" => rgb <= "101111";
					when "100011101111101" => rgb <= "101111";
					when "100011101111110" => rgb <= "101111";
					when "100011101111111" => rgb <= "101111";
					when "100011110000000" => rgb <= "101111";
					when "100011110000001" => rgb <= "101111";
					when "100011110000010" => rgb <= "101111";
					when "100011110000011" => rgb <= "101111";
					when "100011110000100" => rgb <= "101111";
					when "100011110000101" => rgb <= "101111";
					when "100011110000110" => rgb <= "101111";
					when "100011110000111" => rgb <= "101111";
					when "100011110001000" => rgb <= "101111";
					when "100011110001001" => rgb <= "101111";
					when "100011110001010" => rgb <= "101111";
					when "100011110001011" => rgb <= "101111";
					when "100011110001100" => rgb <= "101111";
					when "100011110001101" => rgb <= "101111";
					when "100011110001110" => rgb <= "101111";
					when "100011110001111" => rgb <= "101111";
					when "100011110010000" => rgb <= "101111";
					when "100011110010001" => rgb <= "101111";
					when "100011110010010" => rgb <= "101111";
					when "100011110010011" => rgb <= "101111";
					when "100011110010100" => rgb <= "101111";
					when "100011110010101" => rgb <= "101111";
					when "100011110010110" => rgb <= "101111";
					when "100011110010111" => rgb <= "101111";
					when "100011110011000" => rgb <= "101111";
					when "100011110011001" => rgb <= "101111";
					when "100011110011010" => rgb <= "101111";
					when "100011110011011" => rgb <= "101111";
					when "100011110011100" => rgb <= "101111";
					when "100011110011101" => rgb <= "101111";
					when "100011110011110" => rgb <= "101111";
					when "100011110011111" => rgb <= "101111";
					when "100100000000000" => rgb <= "101111";
					when "100100000000001" => rgb <= "101111";
					when "100100000000010" => rgb <= "101111";
					when "100100000000011" => rgb <= "101111";
					when "100100000000100" => rgb <= "101111";
					when "100100000000101" => rgb <= "101111";
					when "100100000000110" => rgb <= "101111";
					when "100100000000111" => rgb <= "101111";
					when "100100000001000" => rgb <= "101111";
					when "100100000001001" => rgb <= "101111";
					when "100100000001010" => rgb <= "101111";
					when "100100000001011" => rgb <= "101111";
					when "100100000001100" => rgb <= "101111";
					when "100100000001101" => rgb <= "101111";
					when "100100000001110" => rgb <= "101111";
					when "100100000001111" => rgb <= "101111";
					when "100100000010000" => rgb <= "101111";
					when "100100000010001" => rgb <= "101111";
					when "100100000010010" => rgb <= "101111";
					when "100100000010011" => rgb <= "101111";
					when "100100000010100" => rgb <= "101111";
					when "100100000010101" => rgb <= "101111";
					when "100100000010110" => rgb <= "101111";
					when "100100000010111" => rgb <= "101111";
					when "100100000011000" => rgb <= "101111";
					when "100100000011001" => rgb <= "101111";
					when "100100000011010" => rgb <= "101111";
					when "100100000011011" => rgb <= "101111";
					when "100100000011100" => rgb <= "101111";
					when "100100000011101" => rgb <= "101111";
					when "100100000011110" => rgb <= "101111";
					when "100100000011111" => rgb <= "101111";
					when "100100000100000" => rgb <= "000000";
					when "100100000100001" => rgb <= "000000";
					when "100100000100010" => rgb <= "100100";
					when "100100000100011" => rgb <= "100100";
					when "100100000100100" => rgb <= "100100";
					when "100100000100101" => rgb <= "100100";
					when "100100000100110" => rgb <= "000000";
					when "100100000100111" => rgb <= "000000";
					when "100100000101000" => rgb <= "000000";
					when "100100000101001" => rgb <= "000000";
					when "100100000101010" => rgb <= "000000";
					when "100100000101011" => rgb <= "000000";
					when "100100000101100" => rgb <= "100100";
					when "100100000101101" => rgb <= "100100";
					when "100100000101110" => rgb <= "000000";
					when "100100000101111" => rgb <= "000000";
					when "100100000110000" => rgb <= "000000";
					when "100100000110001" => rgb <= "000000";
					when "100100000110010" => rgb <= "000000";
					when "100100000110011" => rgb <= "000000";
					when "100100000110100" => rgb <= "000000";
					when "100100000110101" => rgb <= "000000";
					when "100100000110110" => rgb <= "101111";
					when "100100000110111" => rgb <= "101111";
					when "100100000111000" => rgb <= "101111";
					when "100100000111001" => rgb <= "101111";
					when "100100000111010" => rgb <= "101111";
					when "100100000111011" => rgb <= "101111";
					when "100100000111100" => rgb <= "101111";
					when "100100000111101" => rgb <= "101111";
					when "100100000111110" => rgb <= "101111";
					when "100100000111111" => rgb <= "101111";
					when "100100001000000" => rgb <= "101111";
					when "100100001000001" => rgb <= "101111";
					when "100100001000010" => rgb <= "101111";
					when "100100001000011" => rgb <= "101111";
					when "100100001000100" => rgb <= "101111";
					when "100100001000101" => rgb <= "101111";
					when "100100001000110" => rgb <= "101111";
					when "100100001000111" => rgb <= "101111";
					when "100100001001000" => rgb <= "101111";
					when "100100001001001" => rgb <= "101111";
					when "100100001001010" => rgb <= "101111";
					when "100100001001011" => rgb <= "101111";
					when "100100001001100" => rgb <= "101111";
					when "100100001001101" => rgb <= "101111";
					when "100100001001110" => rgb <= "101111";
					when "100100001001111" => rgb <= "101111";
					when "100100001010000" => rgb <= "101111";
					when "100100001010001" => rgb <= "101111";
					when "100100001010010" => rgb <= "101111";
					when "100100001010011" => rgb <= "101111";
					when "100100001010100" => rgb <= "101111";
					when "100100001010101" => rgb <= "101111";
					when "100100001010110" => rgb <= "101111";
					when "100100001010111" => rgb <= "101111";
					when "100100001011000" => rgb <= "101111";
					when "100100001011001" => rgb <= "101111";
					when "100100001011010" => rgb <= "101111";
					when "100100001011011" => rgb <= "101111";
					when "100100001011100" => rgb <= "101111";
					when "100100001011101" => rgb <= "101111";
					when "100100001011110" => rgb <= "101111";
					when "100100001011111" => rgb <= "101111";
					when "100100001100000" => rgb <= "101111";
					when "100100001100001" => rgb <= "101111";
					when "100100001100010" => rgb <= "101111";
					when "100100001100011" => rgb <= "101111";
					when "100100001100100" => rgb <= "101111";
					when "100100001100101" => rgb <= "101111";
					when "100100001100110" => rgb <= "101111";
					when "100100001100111" => rgb <= "101111";
					when "100100001101000" => rgb <= "101111";
					when "100100001101001" => rgb <= "101111";
					when "100100001101010" => rgb <= "101111";
					when "100100001101011" => rgb <= "101111";
					when "100100001101100" => rgb <= "101111";
					when "100100001101101" => rgb <= "101111";
					when "100100001101110" => rgb <= "101111";
					when "100100001101111" => rgb <= "101111";
					when "100100001110000" => rgb <= "101111";
					when "100100001110001" => rgb <= "101111";
					when "100100001110010" => rgb <= "101111";
					when "100100001110011" => rgb <= "101111";
					when "100100001110100" => rgb <= "101111";
					when "100100001110101" => rgb <= "101111";
					when "100100001110110" => rgb <= "101111";
					when "100100001110111" => rgb <= "101111";
					when "100100001111000" => rgb <= "101111";
					when "100100001111001" => rgb <= "101111";
					when "100100001111010" => rgb <= "101111";
					when "100100001111011" => rgb <= "101111";
					when "100100001111100" => rgb <= "101111";
					when "100100001111101" => rgb <= "101111";
					when "100100001111110" => rgb <= "101111";
					when "100100001111111" => rgb <= "101111";
					when "100100010000000" => rgb <= "101111";
					when "100100010000001" => rgb <= "101111";
					when "100100010000010" => rgb <= "101111";
					when "100100010000011" => rgb <= "101111";
					when "100100010000100" => rgb <= "101111";
					when "100100010000101" => rgb <= "101111";
					when "100100010000110" => rgb <= "101111";
					when "100100010000111" => rgb <= "101111";
					when "100100010001000" => rgb <= "101111";
					when "100100010001001" => rgb <= "101111";
					when "100100010001010" => rgb <= "101111";
					when "100100010001011" => rgb <= "101111";
					when "100100010001100" => rgb <= "101111";
					when "100100010001101" => rgb <= "101111";
					when "100100010001110" => rgb <= "101111";
					when "100100010001111" => rgb <= "101111";
					when "100100010010000" => rgb <= "101111";
					when "100100010010001" => rgb <= "101111";
					when "100100010010010" => rgb <= "101111";
					when "100100010010011" => rgb <= "101111";
					when "100100010010100" => rgb <= "101111";
					when "100100010010101" => rgb <= "101111";
					when "100100010010110" => rgb <= "101111";
					when "100100010010111" => rgb <= "101111";
					when "100100010011000" => rgb <= "101111";
					when "100100010011001" => rgb <= "101111";
					when "100100010011010" => rgb <= "101111";
					when "100100010011011" => rgb <= "101111";
					when "100100010011100" => rgb <= "101111";
					when "100100010011101" => rgb <= "101111";
					when "100100010011110" => rgb <= "101111";
					when "100100010011111" => rgb <= "101111";
					when "100100100000000" => rgb <= "101111";
					when "100100100000001" => rgb <= "101111";
					when "100100100000010" => rgb <= "101111";
					when "100100100000011" => rgb <= "101111";
					when "100100100000100" => rgb <= "101111";
					when "100100100000101" => rgb <= "101111";
					when "100100100000110" => rgb <= "101111";
					when "100100100000111" => rgb <= "101111";
					when "100100100001000" => rgb <= "101111";
					when "100100100001001" => rgb <= "101111";
					when "100100100001010" => rgb <= "101111";
					when "100100100001011" => rgb <= "101111";
					when "100100100001100" => rgb <= "101111";
					when "100100100001101" => rgb <= "101111";
					when "100100100001110" => rgb <= "101111";
					when "100100100001111" => rgb <= "101111";
					when "100100100010000" => rgb <= "101111";
					when "100100100010001" => rgb <= "101111";
					when "100100100010010" => rgb <= "101111";
					when "100100100010011" => rgb <= "101111";
					when "100100100010100" => rgb <= "101111";
					when "100100100010101" => rgb <= "101111";
					when "100100100010110" => rgb <= "101111";
					when "100100100010111" => rgb <= "101111";
					when "100100100011000" => rgb <= "101111";
					when "100100100011001" => rgb <= "101111";
					when "100100100011010" => rgb <= "101111";
					when "100100100011011" => rgb <= "101111";
					when "100100100011100" => rgb <= "101111";
					when "100100100011101" => rgb <= "101111";
					when "100100100011110" => rgb <= "101111";
					when "100100100011111" => rgb <= "101111";
					when "100100100100000" => rgb <= "000000";
					when "100100100100001" => rgb <= "000000";
					when "100100100100010" => rgb <= "100100";
					when "100100100100011" => rgb <= "100100";
					when "100100100100100" => rgb <= "100100";
					when "100100100100101" => rgb <= "100100";
					when "100100100100110" => rgb <= "000000";
					when "100100100100111" => rgb <= "000000";
					when "100100100101000" => rgb <= "000000";
					when "100100100101001" => rgb <= "000000";
					when "100100100101010" => rgb <= "000000";
					when "100100100101011" => rgb <= "000000";
					when "100100100101100" => rgb <= "100100";
					when "100100100101101" => rgb <= "100100";
					when "100100100101110" => rgb <= "000000";
					when "100100100101111" => rgb <= "000000";
					when "100100100110000" => rgb <= "000000";
					when "100100100110001" => rgb <= "000000";
					when "100100100110010" => rgb <= "000000";
					when "100100100110011" => rgb <= "000000";
					when "100100100110100" => rgb <= "000000";
					when "100100100110101" => rgb <= "000000";
					when "100100100110110" => rgb <= "101111";
					when "100100100110111" => rgb <= "101111";
					when "100100100111000" => rgb <= "101111";
					when "100100100111001" => rgb <= "101111";
					when "100100100111010" => rgb <= "101111";
					when "100100100111011" => rgb <= "101111";
					when "100100100111100" => rgb <= "101111";
					when "100100100111101" => rgb <= "101111";
					when "100100100111110" => rgb <= "101111";
					when "100100100111111" => rgb <= "101111";
					when "100100101000000" => rgb <= "101111";
					when "100100101000001" => rgb <= "101111";
					when "100100101000010" => rgb <= "101111";
					when "100100101000011" => rgb <= "101111";
					when "100100101000100" => rgb <= "101111";
					when "100100101000101" => rgb <= "101111";
					when "100100101000110" => rgb <= "101111";
					when "100100101000111" => rgb <= "101111";
					when "100100101001000" => rgb <= "101111";
					when "100100101001001" => rgb <= "101111";
					when "100100101001010" => rgb <= "101111";
					when "100100101001011" => rgb <= "101111";
					when "100100101001100" => rgb <= "101111";
					when "100100101001101" => rgb <= "101111";
					when "100100101001110" => rgb <= "101111";
					when "100100101001111" => rgb <= "101111";
					when "100100101010000" => rgb <= "101111";
					when "100100101010001" => rgb <= "101111";
					when "100100101010010" => rgb <= "101111";
					when "100100101010011" => rgb <= "101111";
					when "100100101010100" => rgb <= "101111";
					when "100100101010101" => rgb <= "101111";
					when "100100101010110" => rgb <= "101111";
					when "100100101010111" => rgb <= "101111";
					when "100100101011000" => rgb <= "101111";
					when "100100101011001" => rgb <= "101111";
					when "100100101011010" => rgb <= "101111";
					when "100100101011011" => rgb <= "101111";
					when "100100101011100" => rgb <= "101111";
					when "100100101011101" => rgb <= "101111";
					when "100100101011110" => rgb <= "101111";
					when "100100101011111" => rgb <= "101111";
					when "100100101100000" => rgb <= "101111";
					when "100100101100001" => rgb <= "101111";
					when "100100101100010" => rgb <= "101111";
					when "100100101100011" => rgb <= "101111";
					when "100100101100100" => rgb <= "101111";
					when "100100101100101" => rgb <= "101111";
					when "100100101100110" => rgb <= "101111";
					when "100100101100111" => rgb <= "101111";
					when "100100101101000" => rgb <= "101111";
					when "100100101101001" => rgb <= "101111";
					when "100100101101010" => rgb <= "101111";
					when "100100101101011" => rgb <= "101111";
					when "100100101101100" => rgb <= "101111";
					when "100100101101101" => rgb <= "101111";
					when "100100101101110" => rgb <= "101111";
					when "100100101101111" => rgb <= "101111";
					when "100100101110000" => rgb <= "101111";
					when "100100101110001" => rgb <= "101111";
					when "100100101110010" => rgb <= "101111";
					when "100100101110011" => rgb <= "101111";
					when "100100101110100" => rgb <= "101111";
					when "100100101110101" => rgb <= "101111";
					when "100100101110110" => rgb <= "101111";
					when "100100101110111" => rgb <= "101111";
					when "100100101111000" => rgb <= "101111";
					when "100100101111001" => rgb <= "101111";
					when "100100101111010" => rgb <= "101111";
					when "100100101111011" => rgb <= "101111";
					when "100100101111100" => rgb <= "101111";
					when "100100101111101" => rgb <= "101111";
					when "100100101111110" => rgb <= "101111";
					when "100100101111111" => rgb <= "101111";
					when "100100110000000" => rgb <= "101111";
					when "100100110000001" => rgb <= "101111";
					when "100100110000010" => rgb <= "101111";
					when "100100110000011" => rgb <= "101111";
					when "100100110000100" => rgb <= "101111";
					when "100100110000101" => rgb <= "101111";
					when "100100110000110" => rgb <= "101111";
					when "100100110000111" => rgb <= "101111";
					when "100100110001000" => rgb <= "101111";
					when "100100110001001" => rgb <= "101111";
					when "100100110001010" => rgb <= "101111";
					when "100100110001011" => rgb <= "101111";
					when "100100110001100" => rgb <= "101111";
					when "100100110001101" => rgb <= "101111";
					when "100100110001110" => rgb <= "101111";
					when "100100110001111" => rgb <= "101111";
					when "100100110010000" => rgb <= "101111";
					when "100100110010001" => rgb <= "101111";
					when "100100110010010" => rgb <= "101111";
					when "100100110010011" => rgb <= "101111";
					when "100100110010100" => rgb <= "101111";
					when "100100110010101" => rgb <= "101111";
					when "100100110010110" => rgb <= "101111";
					when "100100110010111" => rgb <= "101111";
					when "100100110011000" => rgb <= "101111";
					when "100100110011001" => rgb <= "101111";
					when "100100110011010" => rgb <= "101111";
					when "100100110011011" => rgb <= "101111";
					when "100100110011100" => rgb <= "101111";
					when "100100110011101" => rgb <= "101111";
					when "100100110011110" => rgb <= "101111";
					when "100100110011111" => rgb <= "101111";
					when "100101000000000" => rgb <= "101111";
					when "100101000000001" => rgb <= "101111";
					when "100101000000010" => rgb <= "101111";
					when "100101000000011" => rgb <= "101111";
					when "100101000000100" => rgb <= "101111";
					when "100101000000101" => rgb <= "101111";
					when "100101000000110" => rgb <= "101111";
					when "100101000000111" => rgb <= "101111";
					when "100101000001000" => rgb <= "101111";
					when "100101000001001" => rgb <= "101111";
					when "100101000001010" => rgb <= "101111";
					when "100101000001011" => rgb <= "101111";
					when "100101000001100" => rgb <= "101111";
					when "100101000001101" => rgb <= "101111";
					when "100101000001110" => rgb <= "101111";
					when "100101000001111" => rgb <= "101111";
					when "100101000010000" => rgb <= "101111";
					when "100101000010001" => rgb <= "101111";
					when "100101000010010" => rgb <= "101111";
					when "100101000010011" => rgb <= "101111";
					when "100101000010100" => rgb <= "101111";
					when "100101000010101" => rgb <= "101111";
					when "100101000010110" => rgb <= "101111";
					when "100101000010111" => rgb <= "101111";
					when "100101000011000" => rgb <= "101111";
					when "100101000011001" => rgb <= "101111";
					when "100101000011010" => rgb <= "101111";
					when "100101000011011" => rgb <= "101111";
					when "100101000011100" => rgb <= "101111";
					when "100101000011101" => rgb <= "101111";
					when "100101000011110" => rgb <= "101111";
					when "100101000011111" => rgb <= "101111";
					when "100101000100000" => rgb <= "000000";
					when "100101000100001" => rgb <= "000000";
					when "100101000100010" => rgb <= "100100";
					when "100101000100011" => rgb <= "100100";
					when "100101000100100" => rgb <= "100100";
					when "100101000100101" => rgb <= "100100";
					when "100101000100110" => rgb <= "000000";
					when "100101000100111" => rgb <= "000000";
					when "100101000101000" => rgb <= "000000";
					when "100101000101001" => rgb <= "000000";
					when "100101000101010" => rgb <= "000000";
					when "100101000101011" => rgb <= "000000";
					when "100101000101100" => rgb <= "100100";
					when "100101000101101" => rgb <= "100100";
					when "100101000101110" => rgb <= "000000";
					when "100101000101111" => rgb <= "000000";
					when "100101000110000" => rgb <= "000000";
					when "100101000110001" => rgb <= "000000";
					when "100101000110010" => rgb <= "000000";
					when "100101000110011" => rgb <= "000000";
					when "100101000110100" => rgb <= "000010";
					when "100101000110101" => rgb <= "000010";
					when "100101000110110" => rgb <= "000010";
					when "100101000110111" => rgb <= "000010";
					when "100101000111000" => rgb <= "000010";
					when "100101000111001" => rgb <= "000010";
					when "100101000111010" => rgb <= "000010";
					when "100101000111011" => rgb <= "000010";
					when "100101000111100" => rgb <= "000010";
					when "100101000111101" => rgb <= "000010";
					when "100101000111110" => rgb <= "000010";
					when "100101000111111" => rgb <= "000010";
					when "100101001000000" => rgb <= "000010";
					when "100101001000001" => rgb <= "000010";
					when "100101001000010" => rgb <= "000010";
					when "100101001000011" => rgb <= "000010";
					when "100101001000100" => rgb <= "000010";
					when "100101001000101" => rgb <= "000010";
					when "100101001000110" => rgb <= "000010";
					when "100101001000111" => rgb <= "000010";
					when "100101001001000" => rgb <= "000010";
					when "100101001001001" => rgb <= "000010";
					when "100101001001010" => rgb <= "000010";
					when "100101001001011" => rgb <= "000010";
					when "100101001001100" => rgb <= "000010";
					when "100101001001101" => rgb <= "000010";
					when "100101001001110" => rgb <= "000010";
					when "100101001001111" => rgb <= "000010";
					when "100101001010000" => rgb <= "000010";
					when "100101001010001" => rgb <= "000010";
					when "100101001010010" => rgb <= "000010";
					when "100101001010011" => rgb <= "000010";
					when "100101001010100" => rgb <= "000010";
					when "100101001010101" => rgb <= "000010";
					when "100101001010110" => rgb <= "000010";
					when "100101001010111" => rgb <= "000010";
					when "100101001011000" => rgb <= "000010";
					when "100101001011001" => rgb <= "000010";
					when "100101001011010" => rgb <= "000010";
					when "100101001011011" => rgb <= "000010";
					when "100101001011100" => rgb <= "000010";
					when "100101001011101" => rgb <= "000010";
					when "100101001011110" => rgb <= "000010";
					when "100101001011111" => rgb <= "000010";
					when "100101001100000" => rgb <= "000010";
					when "100101001100001" => rgb <= "000010";
					when "100101001100010" => rgb <= "000010";
					when "100101001100011" => rgb <= "000010";
					when "100101001100100" => rgb <= "000010";
					when "100101001100101" => rgb <= "000010";
					when "100101001100110" => rgb <= "000010";
					when "100101001100111" => rgb <= "000010";
					when "100101001101000" => rgb <= "000010";
					when "100101001101001" => rgb <= "000010";
					when "100101001101010" => rgb <= "000010";
					when "100101001101011" => rgb <= "000010";
					when "100101001101100" => rgb <= "101111";
					when "100101001101101" => rgb <= "101111";
					when "100101001101110" => rgb <= "101111";
					when "100101001101111" => rgb <= "101111";
					when "100101001110000" => rgb <= "101111";
					when "100101001110001" => rgb <= "101111";
					when "100101001110010" => rgb <= "101111";
					when "100101001110011" => rgb <= "101111";
					when "100101001110100" => rgb <= "101111";
					when "100101001110101" => rgb <= "101111";
					when "100101001110110" => rgb <= "101111";
					when "100101001110111" => rgb <= "101111";
					when "100101001111000" => rgb <= "101111";
					when "100101001111001" => rgb <= "101111";
					when "100101001111010" => rgb <= "101111";
					when "100101001111011" => rgb <= "101111";
					when "100101001111100" => rgb <= "101111";
					when "100101001111101" => rgb <= "101111";
					when "100101001111110" => rgb <= "101111";
					when "100101001111111" => rgb <= "101111";
					when "100101010000000" => rgb <= "101111";
					when "100101010000001" => rgb <= "101111";
					when "100101010000010" => rgb <= "101111";
					when "100101010000011" => rgb <= "101111";
					when "100101010000100" => rgb <= "101111";
					when "100101010000101" => rgb <= "101111";
					when "100101010000110" => rgb <= "101111";
					when "100101010000111" => rgb <= "101111";
					when "100101010001000" => rgb <= "101111";
					when "100101010001001" => rgb <= "101111";
					when "100101010001010" => rgb <= "101111";
					when "100101010001011" => rgb <= "101111";
					when "100101010001100" => rgb <= "101111";
					when "100101010001101" => rgb <= "101111";
					when "100101010001110" => rgb <= "101111";
					when "100101010001111" => rgb <= "101111";
					when "100101010010000" => rgb <= "101111";
					when "100101010010001" => rgb <= "101111";
					when "100101010010010" => rgb <= "101111";
					when "100101010010011" => rgb <= "101111";
					when "100101010010100" => rgb <= "101111";
					when "100101010010101" => rgb <= "101111";
					when "100101010010110" => rgb <= "101111";
					when "100101010010111" => rgb <= "101111";
					when "100101010011000" => rgb <= "101111";
					when "100101010011001" => rgb <= "101111";
					when "100101010011010" => rgb <= "101111";
					when "100101010011011" => rgb <= "101111";
					when "100101010011100" => rgb <= "101111";
					when "100101010011101" => rgb <= "101111";
					when "100101010011110" => rgb <= "101111";
					when "100101010011111" => rgb <= "101111";
					when "100101100000000" => rgb <= "101111";
					when "100101100000001" => rgb <= "101111";
					when "100101100000010" => rgb <= "101111";
					when "100101100000011" => rgb <= "101111";
					when "100101100000100" => rgb <= "101111";
					when "100101100000101" => rgb <= "101111";
					when "100101100000110" => rgb <= "101111";
					when "100101100000111" => rgb <= "101111";
					when "100101100001000" => rgb <= "101111";
					when "100101100001001" => rgb <= "101111";
					when "100101100001010" => rgb <= "101111";
					when "100101100001011" => rgb <= "101111";
					when "100101100001100" => rgb <= "101111";
					when "100101100001101" => rgb <= "101111";
					when "100101100001110" => rgb <= "101111";
					when "100101100001111" => rgb <= "101111";
					when "100101100010000" => rgb <= "101111";
					when "100101100010001" => rgb <= "101111";
					when "100101100010010" => rgb <= "101111";
					when "100101100010011" => rgb <= "101111";
					when "100101100010100" => rgb <= "101111";
					when "100101100010101" => rgb <= "101111";
					when "100101100010110" => rgb <= "101111";
					when "100101100010111" => rgb <= "101111";
					when "100101100011000" => rgb <= "101111";
					when "100101100011001" => rgb <= "101111";
					when "100101100011010" => rgb <= "101111";
					when "100101100011011" => rgb <= "101111";
					when "100101100011100" => rgb <= "101111";
					when "100101100011101" => rgb <= "101111";
					when "100101100011110" => rgb <= "101111";
					when "100101100011111" => rgb <= "101111";
					when "100101100100000" => rgb <= "000000";
					when "100101100100001" => rgb <= "000000";
					when "100101100100010" => rgb <= "100100";
					when "100101100100011" => rgb <= "100100";
					when "100101100100100" => rgb <= "100100";
					when "100101100100101" => rgb <= "100100";
					when "100101100100110" => rgb <= "000000";
					when "100101100100111" => rgb <= "000000";
					when "100101100101000" => rgb <= "000000";
					when "100101100101001" => rgb <= "000000";
					when "100101100101010" => rgb <= "000000";
					when "100101100101011" => rgb <= "000000";
					when "100101100101100" => rgb <= "100100";
					when "100101100101101" => rgb <= "100100";
					when "100101100101110" => rgb <= "000000";
					when "100101100101111" => rgb <= "000000";
					when "100101100110000" => rgb <= "000000";
					when "100101100110001" => rgb <= "000000";
					when "100101100110010" => rgb <= "000000";
					when "100101100110011" => rgb <= "000000";
					when "100101100110100" => rgb <= "000010";
					when "100101100110101" => rgb <= "000010";
					when "100101100110110" => rgb <= "000010";
					when "100101100110111" => rgb <= "000010";
					when "100101100111000" => rgb <= "000010";
					when "100101100111001" => rgb <= "000010";
					when "100101100111010" => rgb <= "000010";
					when "100101100111011" => rgb <= "000010";
					when "100101100111100" => rgb <= "000010";
					when "100101100111101" => rgb <= "000010";
					when "100101100111110" => rgb <= "000010";
					when "100101100111111" => rgb <= "000010";
					when "100101101000000" => rgb <= "000010";
					when "100101101000001" => rgb <= "000010";
					when "100101101000010" => rgb <= "000010";
					when "100101101000011" => rgb <= "000010";
					when "100101101000100" => rgb <= "000010";
					when "100101101000101" => rgb <= "000010";
					when "100101101000110" => rgb <= "000010";
					when "100101101000111" => rgb <= "000010";
					when "100101101001000" => rgb <= "000010";
					when "100101101001001" => rgb <= "000010";
					when "100101101001010" => rgb <= "000010";
					when "100101101001011" => rgb <= "000010";
					when "100101101001100" => rgb <= "000010";
					when "100101101001101" => rgb <= "000010";
					when "100101101001110" => rgb <= "000010";
					when "100101101001111" => rgb <= "000010";
					when "100101101010000" => rgb <= "000010";
					when "100101101010001" => rgb <= "000010";
					when "100101101010010" => rgb <= "000010";
					when "100101101010011" => rgb <= "000010";
					when "100101101010100" => rgb <= "000010";
					when "100101101010101" => rgb <= "000010";
					when "100101101010110" => rgb <= "000010";
					when "100101101010111" => rgb <= "000010";
					when "100101101011000" => rgb <= "000010";
					when "100101101011001" => rgb <= "000010";
					when "100101101011010" => rgb <= "000010";
					when "100101101011011" => rgb <= "000010";
					when "100101101011100" => rgb <= "000010";
					when "100101101011101" => rgb <= "000010";
					when "100101101011110" => rgb <= "000010";
					when "100101101011111" => rgb <= "000010";
					when "100101101100000" => rgb <= "000010";
					when "100101101100001" => rgb <= "000010";
					when "100101101100010" => rgb <= "000010";
					when "100101101100011" => rgb <= "000010";
					when "100101101100100" => rgb <= "000010";
					when "100101101100101" => rgb <= "000010";
					when "100101101100110" => rgb <= "000010";
					when "100101101100111" => rgb <= "000010";
					when "100101101101000" => rgb <= "000010";
					when "100101101101001" => rgb <= "000010";
					when "100101101101010" => rgb <= "000010";
					when "100101101101011" => rgb <= "000010";
					when "100101101101100" => rgb <= "101111";
					when "100101101101101" => rgb <= "101111";
					when "100101101101110" => rgb <= "101111";
					when "100101101101111" => rgb <= "101111";
					when "100101101110000" => rgb <= "101111";
					when "100101101110001" => rgb <= "101111";
					when "100101101110010" => rgb <= "101111";
					when "100101101110011" => rgb <= "101111";
					when "100101101110100" => rgb <= "101111";
					when "100101101110101" => rgb <= "101111";
					when "100101101110110" => rgb <= "101111";
					when "100101101110111" => rgb <= "101111";
					when "100101101111000" => rgb <= "101111";
					when "100101101111001" => rgb <= "101111";
					when "100101101111010" => rgb <= "101111";
					when "100101101111011" => rgb <= "101111";
					when "100101101111100" => rgb <= "101111";
					when "100101101111101" => rgb <= "101111";
					when "100101101111110" => rgb <= "101111";
					when "100101101111111" => rgb <= "101111";
					when "100101110000000" => rgb <= "101111";
					when "100101110000001" => rgb <= "101111";
					when "100101110000010" => rgb <= "101111";
					when "100101110000011" => rgb <= "101111";
					when "100101110000100" => rgb <= "101111";
					when "100101110000101" => rgb <= "101111";
					when "100101110000110" => rgb <= "101111";
					when "100101110000111" => rgb <= "101111";
					when "100101110001000" => rgb <= "101111";
					when "100101110001001" => rgb <= "101111";
					when "100101110001010" => rgb <= "101111";
					when "100101110001011" => rgb <= "101111";
					when "100101110001100" => rgb <= "101111";
					when "100101110001101" => rgb <= "101111";
					when "100101110001110" => rgb <= "101111";
					when "100101110001111" => rgb <= "101111";
					when "100101110010000" => rgb <= "101111";
					when "100101110010001" => rgb <= "101111";
					when "100101110010010" => rgb <= "101111";
					when "100101110010011" => rgb <= "101111";
					when "100101110010100" => rgb <= "101111";
					when "100101110010101" => rgb <= "101111";
					when "100101110010110" => rgb <= "101111";
					when "100101110010111" => rgb <= "101111";
					when "100101110011000" => rgb <= "101111";
					when "100101110011001" => rgb <= "101111";
					when "100101110011010" => rgb <= "101111";
					when "100101110011011" => rgb <= "101111";
					when "100101110011100" => rgb <= "101111";
					when "100101110011101" => rgb <= "101111";
					when "100101110011110" => rgb <= "101111";
					when "100101110011111" => rgb <= "101111";
					when "100110000000000" => rgb <= "101111";
					when "100110000000001" => rgb <= "101111";
					when "100110000000010" => rgb <= "101111";
					when "100110000000011" => rgb <= "101111";
					when "100110000000100" => rgb <= "101111";
					when "100110000000101" => rgb <= "101111";
					when "100110000000110" => rgb <= "101111";
					when "100110000000111" => rgb <= "101111";
					when "100110000001000" => rgb <= "101111";
					when "100110000001001" => rgb <= "101111";
					when "100110000001010" => rgb <= "101111";
					when "100110000001011" => rgb <= "101111";
					when "100110000001100" => rgb <= "101111";
					when "100110000001101" => rgb <= "101111";
					when "100110000001110" => rgb <= "101111";
					when "100110000001111" => rgb <= "101111";
					when "100110000010000" => rgb <= "101111";
					when "100110000010001" => rgb <= "101111";
					when "100110000010010" => rgb <= "101111";
					when "100110000010011" => rgb <= "101111";
					when "100110000010100" => rgb <= "101111";
					when "100110000010101" => rgb <= "101111";
					when "100110000010110" => rgb <= "101111";
					when "100110000010111" => rgb <= "101111";
					when "100110000011000" => rgb <= "101111";
					when "100110000011001" => rgb <= "101111";
					when "100110000011010" => rgb <= "101111";
					when "100110000011011" => rgb <= "101111";
					when "100110000011100" => rgb <= "101111";
					when "100110000011101" => rgb <= "101111";
					when "100110000011110" => rgb <= "101111";
					when "100110000011111" => rgb <= "101111";
					when "100110000100000" => rgb <= "000000";
					when "100110000100001" => rgb <= "000000";
					when "100110000100010" => rgb <= "100100";
					when "100110000100011" => rgb <= "100100";
					when "100110000100100" => rgb <= "100100";
					when "100110000100101" => rgb <= "100100";
					when "100110000100110" => rgb <= "100100";
					when "100110000100111" => rgb <= "100100";
					when "100110000101000" => rgb <= "000000";
					when "100110000101001" => rgb <= "000000";
					when "100110000101010" => rgb <= "100100";
					when "100110000101011" => rgb <= "100100";
					when "100110000101100" => rgb <= "100100";
					when "100110000101101" => rgb <= "100100";
					when "100110000101110" => rgb <= "100100";
					when "100110000101111" => rgb <= "100100";
					when "100110000110000" => rgb <= "000000";
					when "100110000110001" => rgb <= "000000";
					when "100110000110010" => rgb <= "010000";
					when "100110000110011" => rgb <= "010000";
					when "100110000110100" => rgb <= "000011";
					when "100110000110101" => rgb <= "000011";
					when "100110000110110" => rgb <= "000011";
					when "100110000110111" => rgb <= "000011";
					when "100110000111000" => rgb <= "000011";
					when "100110000111001" => rgb <= "000011";
					when "100110000111010" => rgb <= "000011";
					when "100110000111011" => rgb <= "000011";
					when "100110000111100" => rgb <= "000011";
					when "100110000111101" => rgb <= "000011";
					when "100110000111110" => rgb <= "101111";
					when "100110000111111" => rgb <= "000011";
					when "100110001000000" => rgb <= "000011";
					when "100110001000001" => rgb <= "000011";
					when "100110001000010" => rgb <= "000011";
					when "100110001000011" => rgb <= "000011";
					when "100110001000100" => rgb <= "000011";
					when "100110001000101" => rgb <= "000011";
					when "100110001000110" => rgb <= "000011";
					when "100110001000111" => rgb <= "000011";
					when "100110001001000" => rgb <= "000011";
					when "100110001001001" => rgb <= "000011";
					when "100110001001010" => rgb <= "000011";
					when "100110001001011" => rgb <= "000011";
					when "100110001001100" => rgb <= "000011";
					when "100110001001101" => rgb <= "000011";
					when "100110001001110" => rgb <= "000011";
					when "100110001001111" => rgb <= "000011";
					when "100110001010000" => rgb <= "000011";
					when "100110001010001" => rgb <= "000011";
					when "100110001010010" => rgb <= "000011";
					when "100110001010011" => rgb <= "000011";
					when "100110001010100" => rgb <= "101111";
					when "100110001010101" => rgb <= "000011";
					when "100110001010110" => rgb <= "000011";
					when "100110001010111" => rgb <= "000011";
					when "100110001011000" => rgb <= "000011";
					when "100110001011001" => rgb <= "000011";
					when "100110001011010" => rgb <= "000011";
					when "100110001011011" => rgb <= "000011";
					when "100110001011100" => rgb <= "000011";
					when "100110001011101" => rgb <= "000011";
					when "100110001011110" => rgb <= "000011";
					when "100110001011111" => rgb <= "000011";
					when "100110001100000" => rgb <= "000011";
					when "100110001100001" => rgb <= "000011";
					when "100110001100010" => rgb <= "000011";
					when "100110001100011" => rgb <= "000011";
					when "100110001100100" => rgb <= "000011";
					when "100110001100101" => rgb <= "000011";
					when "100110001100110" => rgb <= "000011";
					when "100110001100111" => rgb <= "000011";
					when "100110001101000" => rgb <= "000011";
					when "100110001101001" => rgb <= "000011";
					when "100110001101010" => rgb <= "000011";
					when "100110001101011" => rgb <= "000011";
					when "100110001101100" => rgb <= "101111";
					when "100110001101101" => rgb <= "101111";
					when "100110001101110" => rgb <= "101111";
					when "100110001101111" => rgb <= "101111";
					when "100110001110000" => rgb <= "101111";
					when "100110001110001" => rgb <= "101111";
					when "100110001110010" => rgb <= "101111";
					when "100110001110011" => rgb <= "101111";
					when "100110001110100" => rgb <= "101111";
					when "100110001110101" => rgb <= "101111";
					when "100110001110110" => rgb <= "101111";
					when "100110001110111" => rgb <= "101111";
					when "100110001111000" => rgb <= "101111";
					when "100110001111001" => rgb <= "101111";
					when "100110001111010" => rgb <= "101111";
					when "100110001111011" => rgb <= "101111";
					when "100110001111100" => rgb <= "101111";
					when "100110001111101" => rgb <= "101111";
					when "100110001111110" => rgb <= "101111";
					when "100110001111111" => rgb <= "101111";
					when "100110010000000" => rgb <= "101111";
					when "100110010000001" => rgb <= "101111";
					when "100110010000010" => rgb <= "101111";
					when "100110010000011" => rgb <= "101111";
					when "100110010000100" => rgb <= "101111";
					when "100110010000101" => rgb <= "101111";
					when "100110010000110" => rgb <= "101111";
					when "100110010000111" => rgb <= "101111";
					when "100110010001000" => rgb <= "101111";
					when "100110010001001" => rgb <= "101111";
					when "100110010001010" => rgb <= "101111";
					when "100110010001011" => rgb <= "101111";
					when "100110010001100" => rgb <= "101111";
					when "100110010001101" => rgb <= "101111";
					when "100110010001110" => rgb <= "101111";
					when "100110010001111" => rgb <= "101111";
					when "100110010010000" => rgb <= "101111";
					when "100110010010001" => rgb <= "101111";
					when "100110010010010" => rgb <= "101111";
					when "100110010010011" => rgb <= "101111";
					when "100110010010100" => rgb <= "101111";
					when "100110010010101" => rgb <= "101111";
					when "100110010010110" => rgb <= "101111";
					when "100110010010111" => rgb <= "101111";
					when "100110010011000" => rgb <= "101111";
					when "100110010011001" => rgb <= "101111";
					when "100110010011010" => rgb <= "101111";
					when "100110010011011" => rgb <= "101111";
					when "100110010011100" => rgb <= "101111";
					when "100110010011101" => rgb <= "101111";
					when "100110010011110" => rgb <= "101111";
					when "100110010011111" => rgb <= "101111";
					when "100110100000000" => rgb <= "101111";
					when "100110100000001" => rgb <= "101111";
					when "100110100000010" => rgb <= "101111";
					when "100110100000011" => rgb <= "101111";
					when "100110100000100" => rgb <= "101111";
					when "100110100000101" => rgb <= "101111";
					when "100110100000110" => rgb <= "101111";
					when "100110100000111" => rgb <= "101111";
					when "100110100001000" => rgb <= "101111";
					when "100110100001001" => rgb <= "101111";
					when "100110100001010" => rgb <= "101111";
					when "100110100001011" => rgb <= "101111";
					when "100110100001100" => rgb <= "101111";
					when "100110100001101" => rgb <= "101111";
					when "100110100001110" => rgb <= "101111";
					when "100110100001111" => rgb <= "101111";
					when "100110100010000" => rgb <= "101111";
					when "100110100010001" => rgb <= "101111";
					when "100110100010010" => rgb <= "101111";
					when "100110100010011" => rgb <= "101111";
					when "100110100010100" => rgb <= "101111";
					when "100110100010101" => rgb <= "101111";
					when "100110100010110" => rgb <= "101111";
					when "100110100010111" => rgb <= "101111";
					when "100110100011000" => rgb <= "101111";
					when "100110100011001" => rgb <= "101111";
					when "100110100011010" => rgb <= "101111";
					when "100110100011011" => rgb <= "101111";
					when "100110100011100" => rgb <= "101111";
					when "100110100011101" => rgb <= "101111";
					when "100110100011110" => rgb <= "101111";
					when "100110100011111" => rgb <= "101111";
					when "100110100100000" => rgb <= "000000";
					when "100110100100001" => rgb <= "000000";
					when "100110100100010" => rgb <= "100100";
					when "100110100100011" => rgb <= "100100";
					when "100110100100100" => rgb <= "100100";
					when "100110100100101" => rgb <= "100100";
					when "100110100100110" => rgb <= "100100";
					when "100110100100111" => rgb <= "100100";
					when "100110100101000" => rgb <= "000000";
					when "100110100101001" => rgb <= "000000";
					when "100110100101010" => rgb <= "100100";
					when "100110100101011" => rgb <= "100100";
					when "100110100101100" => rgb <= "100100";
					when "100110100101101" => rgb <= "100100";
					when "100110100101110" => rgb <= "100100";
					when "100110100101111" => rgb <= "100100";
					when "100110100110000" => rgb <= "000000";
					when "100110100110001" => rgb <= "000000";
					when "100110100110010" => rgb <= "010000";
					when "100110100110011" => rgb <= "010000";
					when "100110100110100" => rgb <= "000000";
					when "100110100110101" => rgb <= "000000";
					when "100110100110110" => rgb <= "000011";
					when "100110100110111" => rgb <= "000011";
					when "100110100111000" => rgb <= "000011";
					when "100110100111001" => rgb <= "000011";
					when "100110100111010" => rgb <= "000011";
					when "100110100111011" => rgb <= "101111";
					when "100110100111100" => rgb <= "101111";
					when "100110100111101" => rgb <= "101111";
					when "100110100111110" => rgb <= "101111";
					when "100110100111111" => rgb <= "101111";
					when "100110101000000" => rgb <= "101111";
					when "100110101000001" => rgb <= "000011";
					when "100110101000010" => rgb <= "000011";
					when "100110101000011" => rgb <= "000011";
					when "100110101000100" => rgb <= "000011";
					when "100110101000101" => rgb <= "000011";
					when "100110101000110" => rgb <= "000011";
					when "100110101000111" => rgb <= "000011";
					when "100110101001000" => rgb <= "101111";
					when "100110101001001" => rgb <= "000011";
					when "100110101001010" => rgb <= "101111";
					when "100110101001011" => rgb <= "000011";
					when "100110101001100" => rgb <= "000011";
					when "100110101001101" => rgb <= "000011";
					when "100110101001110" => rgb <= "101111";
					when "100110101001111" => rgb <= "000011";
					when "100110101010000" => rgb <= "000011";
					when "100110101010001" => rgb <= "000011";
					when "100110101010010" => rgb <= "000011";
					when "100110101010011" => rgb <= "000011";
					when "100110101010100" => rgb <= "101111";
					when "100110101010101" => rgb <= "101111";
					when "100110101010110" => rgb <= "000011";
					when "100110101010111" => rgb <= "000011";
					when "100110101011000" => rgb <= "000011";
					when "100110101011001" => rgb <= "000011";
					when "100110101011010" => rgb <= "101111";
					when "100110101011011" => rgb <= "101111";
					when "100110101011100" => rgb <= "101111";
					when "100110101011101" => rgb <= "000011";
					when "100110101011110" => rgb <= "101111";
					when "100110101011111" => rgb <= "101111";
					when "100110101100000" => rgb <= "000011";
					when "100110101100001" => rgb <= "000011";
					when "100110101100010" => rgb <= "000011";
					when "100110101100011" => rgb <= "101111";
					when "100110101100100" => rgb <= "000011";
					when "100110101100101" => rgb <= "000011";
					when "100110101100110" => rgb <= "101111";
					when "100110101100111" => rgb <= "000011";
					when "100110101101000" => rgb <= "000011";
					when "100110101101001" => rgb <= "000011";
					when "100110101101010" => rgb <= "101111";
					when "100110101101011" => rgb <= "101111";
					when "100110101101100" => rgb <= "101111";
					when "100110101101101" => rgb <= "101111";
					when "100110101101110" => rgb <= "101111";
					when "100110101101111" => rgb <= "101111";
					when "100110101110000" => rgb <= "101111";
					when "100110101110001" => rgb <= "101111";
					when "100110101110010" => rgb <= "101111";
					when "100110101110011" => rgb <= "101111";
					when "100110101110100" => rgb <= "101111";
					when "100110101110101" => rgb <= "101111";
					when "100110101110110" => rgb <= "101111";
					when "100110101110111" => rgb <= "101111";
					when "100110101111000" => rgb <= "101111";
					when "100110101111001" => rgb <= "101111";
					when "100110101111010" => rgb <= "101111";
					when "100110101111011" => rgb <= "101111";
					when "100110101111100" => rgb <= "101111";
					when "100110101111101" => rgb <= "101111";
					when "100110101111110" => rgb <= "101111";
					when "100110101111111" => rgb <= "101111";
					when "100110110000000" => rgb <= "101111";
					when "100110110000001" => rgb <= "101111";
					when "100110110000010" => rgb <= "101111";
					when "100110110000011" => rgb <= "101111";
					when "100110110000100" => rgb <= "101111";
					when "100110110000101" => rgb <= "101111";
					when "100110110000110" => rgb <= "101111";
					when "100110110000111" => rgb <= "101111";
					when "100110110001000" => rgb <= "101111";
					when "100110110001001" => rgb <= "101111";
					when "100110110001010" => rgb <= "101111";
					when "100110110001011" => rgb <= "101111";
					when "100110110001100" => rgb <= "101111";
					when "100110110001101" => rgb <= "101111";
					when "100110110001110" => rgb <= "101111";
					when "100110110001111" => rgb <= "101111";
					when "100110110010000" => rgb <= "101111";
					when "100110110010001" => rgb <= "101111";
					when "100110110010010" => rgb <= "101111";
					when "100110110010011" => rgb <= "101111";
					when "100110110010100" => rgb <= "101111";
					when "100110110010101" => rgb <= "101111";
					when "100110110010110" => rgb <= "101111";
					when "100110110010111" => rgb <= "101111";
					when "100110110011000" => rgb <= "101111";
					when "100110110011001" => rgb <= "101111";
					when "100110110011010" => rgb <= "101111";
					when "100110110011011" => rgb <= "101111";
					when "100110110011100" => rgb <= "101111";
					when "100110110011101" => rgb <= "101111";
					when "100110110011110" => rgb <= "101111";
					when "100110110011111" => rgb <= "101111";
					when "100111000000000" => rgb <= "101111";
					when "100111000000001" => rgb <= "101111";
					when "100111000000010" => rgb <= "101111";
					when "100111000000011" => rgb <= "101111";
					when "100111000000100" => rgb <= "101111";
					when "100111000000101" => rgb <= "101111";
					when "100111000000110" => rgb <= "101111";
					when "100111000000111" => rgb <= "101111";
					when "100111000001000" => rgb <= "101111";
					when "100111000001001" => rgb <= "101111";
					when "100111000001010" => rgb <= "101111";
					when "100111000001011" => rgb <= "101111";
					when "100111000001100" => rgb <= "101111";
					when "100111000001101" => rgb <= "101111";
					when "100111000001110" => rgb <= "101111";
					when "100111000001111" => rgb <= "101111";
					when "100111000010000" => rgb <= "101111";
					when "100111000010001" => rgb <= "101111";
					when "100111000010010" => rgb <= "101111";
					when "100111000010011" => rgb <= "101111";
					when "100111000010100" => rgb <= "101111";
					when "100111000010101" => rgb <= "101111";
					when "100111000010110" => rgb <= "101111";
					when "100111000010111" => rgb <= "101111";
					when "100111000011000" => rgb <= "101111";
					when "100111000011001" => rgb <= "101111";
					when "100111000011010" => rgb <= "101111";
					when "100111000011011" => rgb <= "101111";
					when "100111000011100" => rgb <= "101111";
					when "100111000011101" => rgb <= "101111";
					when "100111000011110" => rgb <= "101111";
					when "100111000011111" => rgb <= "101111";
					when "100111000100000" => rgb <= "000000";
					when "100111000100001" => rgb <= "000000";
					when "100111000100010" => rgb <= "100100";
					when "100111000100011" => rgb <= "100100";
					when "100111000100100" => rgb <= "100100";
					when "100111000100101" => rgb <= "100100";
					when "100111000100110" => rgb <= "100100";
					when "100111000100111" => rgb <= "100100";
					when "100111000101000" => rgb <= "100100";
					when "100111000101001" => rgb <= "100100";
					when "100111000101010" => rgb <= "100100";
					when "100111000101011" => rgb <= "100100";
					when "100111000101100" => rgb <= "100100";
					when "100111000101101" => rgb <= "100100";
					when "100111000101110" => rgb <= "100100";
					when "100111000101111" => rgb <= "100100";
					when "100111000110000" => rgb <= "100100";
					when "100111000110001" => rgb <= "100100";
					when "100111000110010" => rgb <= "010000";
					when "100111000110011" => rgb <= "010000";
					when "100111000110100" => rgb <= "000000";
					when "100111000110101" => rgb <= "000000";
					when "100111000110110" => rgb <= "101111";
					when "100111000110111" => rgb <= "101111";
					when "100111000111000" => rgb <= "101111";
					when "100111000111001" => rgb <= "000011";
					when "100111000111010" => rgb <= "101111";
					when "100111000111011" => rgb <= "101111";
					when "100111000111100" => rgb <= "101111";
					when "100111000111101" => rgb <= "101111";
					when "100111000111110" => rgb <= "101111";
					when "100111000111111" => rgb <= "101111";
					when "100111001000000" => rgb <= "101111";
					when "100111001000001" => rgb <= "101111";
					when "100111001000010" => rgb <= "000011";
					when "100111001000011" => rgb <= "101111";
					when "100111001000100" => rgb <= "101111";
					when "100111001000101" => rgb <= "000011";
					when "100111001000110" => rgb <= "000011";
					when "100111001000111" => rgb <= "101111";
					when "100111001001000" => rgb <= "101111";
					when "100111001001001" => rgb <= "101111";
					when "100111001001010" => rgb <= "101111";
					when "100111001001011" => rgb <= "000011";
					when "100111001001100" => rgb <= "000011";
					when "100111001001101" => rgb <= "101111";
					when "100111001001110" => rgb <= "101111";
					when "100111001001111" => rgb <= "101111";
					when "100111001010000" => rgb <= "101111";
					when "100111001010001" => rgb <= "000011";
					when "100111001010010" => rgb <= "101111";
					when "100111001010011" => rgb <= "101111";
					when "100111001010100" => rgb <= "101111";
					when "100111001010101" => rgb <= "101111";
					when "100111001010110" => rgb <= "101111";
					when "100111001010111" => rgb <= "101111";
					when "100111001011000" => rgb <= "000011";
					when "100111001011001" => rgb <= "101111";
					when "100111001011010" => rgb <= "101111";
					when "100111001011011" => rgb <= "101111";
					when "100111001011100" => rgb <= "101111";
					when "100111001011101" => rgb <= "101111";
					when "100111001011110" => rgb <= "101111";
					when "100111001011111" => rgb <= "101111";
					when "100111001100000" => rgb <= "101111";
					when "100111001100001" => rgb <= "101111";
					when "100111001100010" => rgb <= "000011";
					when "100111001100011" => rgb <= "101111";
					when "100111001100100" => rgb <= "000011";
					when "100111001100101" => rgb <= "101111";
					when "100111001100110" => rgb <= "101111";
					when "100111001100111" => rgb <= "101111";
					when "100111001101000" => rgb <= "000011";
					when "100111001101001" => rgb <= "101111";
					when "100111001101010" => rgb <= "101111";
					when "100111001101011" => rgb <= "101111";
					when "100111001101100" => rgb <= "101111";
					when "100111001101101" => rgb <= "101111";
					when "100111001101110" => rgb <= "101111";
					when "100111001101111" => rgb <= "101111";
					when "100111001110000" => rgb <= "101111";
					when "100111001110001" => rgb <= "101111";
					when "100111001110010" => rgb <= "101111";
					when "100111001110011" => rgb <= "101111";
					when "100111001110100" => rgb <= "101111";
					when "100111001110101" => rgb <= "101111";
					when "100111001110110" => rgb <= "101111";
					when "100111001110111" => rgb <= "101111";
					when "100111001111000" => rgb <= "101111";
					when "100111001111001" => rgb <= "101111";
					when "100111001111010" => rgb <= "101111";
					when "100111001111011" => rgb <= "101111";
					when "100111001111100" => rgb <= "101111";
					when "100111001111101" => rgb <= "101111";
					when "100111001111110" => rgb <= "101111";
					when "100111001111111" => rgb <= "101111";
					when "100111010000000" => rgb <= "101111";
					when "100111010000001" => rgb <= "101111";
					when "100111010000010" => rgb <= "101111";
					when "100111010000011" => rgb <= "101111";
					when "100111010000100" => rgb <= "101111";
					when "100111010000101" => rgb <= "101111";
					when "100111010000110" => rgb <= "101111";
					when "100111010000111" => rgb <= "101111";
					when "100111010001000" => rgb <= "101111";
					when "100111010001001" => rgb <= "101111";
					when "100111010001010" => rgb <= "101111";
					when "100111010001011" => rgb <= "101111";
					when "100111010001100" => rgb <= "101111";
					when "100111010001101" => rgb <= "101111";
					when "100111010001110" => rgb <= "101111";
					when "100111010001111" => rgb <= "101111";
					when "100111010010000" => rgb <= "101111";
					when "100111010010001" => rgb <= "101111";
					when "100111010010010" => rgb <= "101111";
					when "100111010010011" => rgb <= "101111";
					when "100111010010100" => rgb <= "101111";
					when "100111010010101" => rgb <= "101111";
					when "100111010010110" => rgb <= "101111";
					when "100111010010111" => rgb <= "101111";
					when "100111010011000" => rgb <= "101111";
					when "100111010011001" => rgb <= "101111";
					when "100111010011010" => rgb <= "101111";
					when "100111010011011" => rgb <= "101111";
					when "100111010011100" => rgb <= "101111";
					when "100111010011101" => rgb <= "101111";
					when "100111010011110" => rgb <= "101111";
					when "100111010011111" => rgb <= "101111";
					when "100111100000000" => rgb <= "101111";
					when "100111100000001" => rgb <= "101111";
					when "100111100000010" => rgb <= "101111";
					when "100111100000011" => rgb <= "101111";
					when "100111100000100" => rgb <= "101111";
					when "100111100000101" => rgb <= "101111";
					when "100111100000110" => rgb <= "101111";
					when "100111100000111" => rgb <= "101111";
					when "100111100001000" => rgb <= "101111";
					when "100111100001001" => rgb <= "101111";
					when "100111100001010" => rgb <= "101111";
					when "100111100001011" => rgb <= "101111";
					when "100111100001100" => rgb <= "101111";
					when "100111100001101" => rgb <= "101111";
					when "100111100001110" => rgb <= "101111";
					when "100111100001111" => rgb <= "101111";
					when "100111100010000" => rgb <= "101111";
					when "100111100010001" => rgb <= "101111";
					when "100111100010010" => rgb <= "101111";
					when "100111100010011" => rgb <= "101111";
					when "100111100010100" => rgb <= "101111";
					when "100111100010101" => rgb <= "101111";
					when "100111100010110" => rgb <= "101111";
					when "100111100010111" => rgb <= "101111";
					when "100111100011000" => rgb <= "101111";
					when "100111100011001" => rgb <= "101111";
					when "100111100011010" => rgb <= "101111";
					when "100111100011011" => rgb <= "101111";
					when "100111100011100" => rgb <= "101111";
					when "100111100011101" => rgb <= "101111";
					when "100111100011110" => rgb <= "101111";
					when "100111100011111" => rgb <= "101111";
					when "100111100100000" => rgb <= "000000";
					when "100111100100001" => rgb <= "000000";
					when "100111100100010" => rgb <= "100100";
					when "100111100100011" => rgb <= "100100";
					when "100111100100100" => rgb <= "100100";
					when "100111100100101" => rgb <= "100100";
					when "100111100100110" => rgb <= "100100";
					when "100111100100111" => rgb <= "100100";
					when "100111100101000" => rgb <= "100100";
					when "100111100101001" => rgb <= "100100";
					when "100111100101010" => rgb <= "100100";
					when "100111100101011" => rgb <= "100100";
					when "100111100101100" => rgb <= "100100";
					when "100111100101101" => rgb <= "100100";
					when "100111100101110" => rgb <= "100100";
					when "100111100101111" => rgb <= "100100";
					when "100111100110000" => rgb <= "100100";
					when "100111100110001" => rgb <= "100100";
					when "100111100110010" => rgb <= "010000";
					when "100111100110011" => rgb <= "010000";
					when "100111100110100" => rgb <= "000000";
					when "100111100110101" => rgb <= "000000";
					when "100111100110110" => rgb <= "101111";
					when "100111100110111" => rgb <= "101111";
					when "100111100111000" => rgb <= "101111";
					when "100111100111001" => rgb <= "101111";
					when "100111100111010" => rgb <= "101111";
					when "100111100111011" => rgb <= "101111";
					when "100111100111100" => rgb <= "101111";
					when "100111100111101" => rgb <= "101111";
					when "100111100111110" => rgb <= "101111";
					when "100111100111111" => rgb <= "101111";
					when "100111101000000" => rgb <= "101111";
					when "100111101000001" => rgb <= "101111";
					when "100111101000010" => rgb <= "101111";
					when "100111101000011" => rgb <= "101111";
					when "100111101000100" => rgb <= "101111";
					when "100111101000101" => rgb <= "101111";
					when "100111101000110" => rgb <= "000011";
					when "100111101000111" => rgb <= "101111";
					when "100111101001000" => rgb <= "101111";
					when "100111101001001" => rgb <= "101111";
					when "100111101001010" => rgb <= "101111";
					when "100111101001011" => rgb <= "000011";
					when "100111101001100" => rgb <= "000011";
					when "100111101001101" => rgb <= "101111";
					when "100111101001110" => rgb <= "101111";
					when "100111101001111" => rgb <= "101111";
					when "100111101010000" => rgb <= "101111";
					when "100111101010001" => rgb <= "101111";
					when "100111101010010" => rgb <= "101111";
					when "100111101010011" => rgb <= "101111";
					when "100111101010100" => rgb <= "101111";
					when "100111101010101" => rgb <= "101111";
					when "100111101010110" => rgb <= "101111";
					when "100111101010111" => rgb <= "101111";
					when "100111101011000" => rgb <= "101111";
					when "100111101011001" => rgb <= "101111";
					when "100111101011010" => rgb <= "101111";
					when "100111101011011" => rgb <= "101111";
					when "100111101011100" => rgb <= "101111";
					when "100111101011101" => rgb <= "101111";
					when "100111101011110" => rgb <= "101111";
					when "100111101011111" => rgb <= "101111";
					when "100111101100000" => rgb <= "101111";
					when "100111101100001" => rgb <= "101111";
					when "100111101100010" => rgb <= "101111";
					when "100111101100011" => rgb <= "101111";
					when "100111101100100" => rgb <= "101111";
					when "100111101100101" => rgb <= "101111";
					when "100111101100110" => rgb <= "101111";
					when "100111101100111" => rgb <= "101111";
					when "100111101101000" => rgb <= "101111";
					when "100111101101001" => rgb <= "101111";
					when "100111101101010" => rgb <= "101111";
					when "100111101101011" => rgb <= "101111";
					when "100111101101100" => rgb <= "101111";
					when "100111101101101" => rgb <= "101111";
					when "100111101101110" => rgb <= "101111";
					when "100111101101111" => rgb <= "101111";
					when "100111101110000" => rgb <= "101111";
					when "100111101110001" => rgb <= "101111";
					when "100111101110010" => rgb <= "101111";
					when "100111101110011" => rgb <= "101111";
					when "100111101110100" => rgb <= "101111";
					when "100111101110101" => rgb <= "101111";
					when "100111101110110" => rgb <= "101111";
					when "100111101110111" => rgb <= "101111";
					when "100111101111000" => rgb <= "101111";
					when "100111101111001" => rgb <= "101111";
					when "100111101111010" => rgb <= "101111";
					when "100111101111011" => rgb <= "101111";
					when "100111101111100" => rgb <= "101111";
					when "100111101111101" => rgb <= "101111";
					when "100111101111110" => rgb <= "101111";
					when "100111101111111" => rgb <= "101111";
					when "100111110000000" => rgb <= "101111";
					when "100111110000001" => rgb <= "101111";
					when "100111110000010" => rgb <= "101111";
					when "100111110000011" => rgb <= "101111";
					when "100111110000100" => rgb <= "101111";
					when "100111110000101" => rgb <= "101111";
					when "100111110000110" => rgb <= "101111";
					when "100111110000111" => rgb <= "101111";
					when "100111110001000" => rgb <= "101111";
					when "100111110001001" => rgb <= "101111";
					when "100111110001010" => rgb <= "101111";
					when "100111110001011" => rgb <= "101111";
					when "100111110001100" => rgb <= "101111";
					when "100111110001101" => rgb <= "101111";
					when "100111110001110" => rgb <= "101111";
					when "100111110001111" => rgb <= "101111";
					when "100111110010000" => rgb <= "101111";
					when "100111110010001" => rgb <= "101111";
					when "100111110010010" => rgb <= "101111";
					when "100111110010011" => rgb <= "101111";
					when "100111110010100" => rgb <= "101111";
					when "100111110010101" => rgb <= "101111";
					when "100111110010110" => rgb <= "101111";
					when "100111110010111" => rgb <= "101111";
					when "100111110011000" => rgb <= "101111";
					when "100111110011001" => rgb <= "101111";
					when "100111110011010" => rgb <= "101111";
					when "100111110011011" => rgb <= "101111";
					when "100111110011100" => rgb <= "101111";
					when "100111110011101" => rgb <= "101111";
					when "100111110011110" => rgb <= "101111";
					when "100111110011111" => rgb <= "101111";
					when "101000000000000" => rgb <= "101111";
					when "101000000000001" => rgb <= "101111";
					when "101000000000010" => rgb <= "101111";
					when "101000000000011" => rgb <= "101111";
					when "101000000000100" => rgb <= "101111";
					when "101000000000101" => rgb <= "101111";
					when "101000000000110" => rgb <= "101111";
					when "101000000000111" => rgb <= "101111";
					when "101000000001000" => rgb <= "101111";
					when "101000000001001" => rgb <= "101111";
					when "101000000001010" => rgb <= "101111";
					when "101000000001011" => rgb <= "101111";
					when "101000000001100" => rgb <= "101111";
					when "101000000001101" => rgb <= "101111";
					when "101000000001110" => rgb <= "101111";
					when "101000000001111" => rgb <= "101111";
					when "101000000010000" => rgb <= "101111";
					when "101000000010001" => rgb <= "101111";
					when "101000000010010" => rgb <= "101111";
					when "101000000010011" => rgb <= "101111";
					when "101000000010100" => rgb <= "101111";
					when "101000000010101" => rgb <= "101111";
					when "101000000010110" => rgb <= "101111";
					when "101000000010111" => rgb <= "101111";
					when "101000000011000" => rgb <= "101111";
					when "101000000011001" => rgb <= "101111";
					when "101000000011010" => rgb <= "101111";
					when "101000000011011" => rgb <= "101111";
					when "101000000011100" => rgb <= "101111";
					when "101000000011101" => rgb <= "101111";
					when "101000000011110" => rgb <= "101111";
					when "101000000011111" => rgb <= "101111";
					when "101000000100000" => rgb <= "000000";
					when "101000000100001" => rgb <= "000000";
					when "101000000100010" => rgb <= "100100";
					when "101000000100011" => rgb <= "100100";
					when "101000000100100" => rgb <= "100100";
					when "101000000100101" => rgb <= "100100";
					when "101000000100110" => rgb <= "100100";
					when "101000000100111" => rgb <= "100100";
					when "101000000101000" => rgb <= "100100";
					when "101000000101001" => rgb <= "100100";
					when "101000000101010" => rgb <= "100100";
					when "101000000101011" => rgb <= "100100";
					when "101000000101100" => rgb <= "000000";
					when "101000000101101" => rgb <= "000000";
					when "101000000101110" => rgb <= "100100";
					when "101000000101111" => rgb <= "100100";
					when "101000000110000" => rgb <= "100100";
					when "101000000110001" => rgb <= "100100";
					when "101000000110010" => rgb <= "010000";
					when "101000000110011" => rgb <= "010000";
					when "101000000110100" => rgb <= "000000";
					when "101000000110101" => rgb <= "000000";
					when "101000000110110" => rgb <= "101111";
					when "101000000110111" => rgb <= "101111";
					when "101000000111000" => rgb <= "101111";
					when "101000000111001" => rgb <= "101111";
					when "101000000111010" => rgb <= "101111";
					when "101000000111011" => rgb <= "101111";
					when "101000000111100" => rgb <= "101111";
					when "101000000111101" => rgb <= "101111";
					when "101000000111110" => rgb <= "101111";
					when "101000000111111" => rgb <= "101111";
					when "101000001000000" => rgb <= "101111";
					when "101000001000001" => rgb <= "101111";
					when "101000001000010" => rgb <= "101111";
					when "101000001000011" => rgb <= "101111";
					when "101000001000100" => rgb <= "101111";
					when "101000001000101" => rgb <= "101111";
					when "101000001000110" => rgb <= "101111";
					when "101000001000111" => rgb <= "101111";
					when "101000001001000" => rgb <= "101111";
					when "101000001001001" => rgb <= "101111";
					when "101000001001010" => rgb <= "101111";
					when "101000001001011" => rgb <= "000011";
					when "101000001001100" => rgb <= "101111";
					when "101000001001101" => rgb <= "101111";
					when "101000001001110" => rgb <= "101111";
					when "101000001001111" => rgb <= "101111";
					when "101000001010000" => rgb <= "101111";
					when "101000001010001" => rgb <= "101111";
					when "101000001010010" => rgb <= "101111";
					when "101000001010011" => rgb <= "101111";
					when "101000001010100" => rgb <= "101111";
					when "101000001010101" => rgb <= "101111";
					when "101000001010110" => rgb <= "101111";
					when "101000001010111" => rgb <= "101111";
					when "101000001011000" => rgb <= "101111";
					when "101000001011001" => rgb <= "101111";
					when "101000001011010" => rgb <= "101111";
					when "101000001011011" => rgb <= "101111";
					when "101000001011100" => rgb <= "101111";
					when "101000001011101" => rgb <= "101111";
					when "101000001011110" => rgb <= "101111";
					when "101000001011111" => rgb <= "101111";
					when "101000001100000" => rgb <= "101111";
					when "101000001100001" => rgb <= "101111";
					when "101000001100010" => rgb <= "101111";
					when "101000001100011" => rgb <= "101111";
					when "101000001100100" => rgb <= "101111";
					when "101000001100101" => rgb <= "101111";
					when "101000001100110" => rgb <= "101111";
					when "101000001100111" => rgb <= "101111";
					when "101000001101000" => rgb <= "101111";
					when "101000001101001" => rgb <= "101111";
					when "101000001101010" => rgb <= "101111";
					when "101000001101011" => rgb <= "101111";
					when "101000001101100" => rgb <= "101111";
					when "101000001101101" => rgb <= "101111";
					when "101000001101110" => rgb <= "101111";
					when "101000001101111" => rgb <= "101111";
					when "101000001110000" => rgb <= "101111";
					when "101000001110001" => rgb <= "101111";
					when "101000001110010" => rgb <= "101111";
					when "101000001110011" => rgb <= "101111";
					when "101000001110100" => rgb <= "101111";
					when "101000001110101" => rgb <= "101111";
					when "101000001110110" => rgb <= "101111";
					when "101000001110111" => rgb <= "101111";
					when "101000001111000" => rgb <= "101111";
					when "101000001111001" => rgb <= "101111";
					when "101000001111010" => rgb <= "101111";
					when "101000001111011" => rgb <= "101111";
					when "101000001111100" => rgb <= "101111";
					when "101000001111101" => rgb <= "101111";
					when "101000001111110" => rgb <= "101111";
					when "101000001111111" => rgb <= "101111";
					when "101000010000000" => rgb <= "101111";
					when "101000010000001" => rgb <= "101111";
					when "101000010000010" => rgb <= "101111";
					when "101000010000011" => rgb <= "101111";
					when "101000010000100" => rgb <= "101111";
					when "101000010000101" => rgb <= "101111";
					when "101000010000110" => rgb <= "101111";
					when "101000010000111" => rgb <= "101111";
					when "101000010001000" => rgb <= "101111";
					when "101000010001001" => rgb <= "101111";
					when "101000010001010" => rgb <= "101111";
					when "101000010001011" => rgb <= "101111";
					when "101000010001100" => rgb <= "101111";
					when "101000010001101" => rgb <= "101111";
					when "101000010001110" => rgb <= "101111";
					when "101000010001111" => rgb <= "101111";
					when "101000010010000" => rgb <= "101111";
					when "101000010010001" => rgb <= "101111";
					when "101000010010010" => rgb <= "101111";
					when "101000010010011" => rgb <= "101111";
					when "101000010010100" => rgb <= "101111";
					when "101000010010101" => rgb <= "101111";
					when "101000010010110" => rgb <= "101111";
					when "101000010010111" => rgb <= "101111";
					when "101000010011000" => rgb <= "101111";
					when "101000010011001" => rgb <= "101111";
					when "101000010011010" => rgb <= "101111";
					when "101000010011011" => rgb <= "101111";
					when "101000010011100" => rgb <= "101111";
					when "101000010011101" => rgb <= "101111";
					when "101000010011110" => rgb <= "101111";
					when "101000010011111" => rgb <= "101111";
					when "101000100000000" => rgb <= "101111";
					when "101000100000001" => rgb <= "101111";
					when "101000100000010" => rgb <= "101111";
					when "101000100000011" => rgb <= "101111";
					when "101000100000100" => rgb <= "101111";
					when "101000100000101" => rgb <= "101111";
					when "101000100000110" => rgb <= "101111";
					when "101000100000111" => rgb <= "101111";
					when "101000100001000" => rgb <= "101111";
					when "101000100001001" => rgb <= "101111";
					when "101000100001010" => rgb <= "101111";
					when "101000100001011" => rgb <= "101111";
					when "101000100001100" => rgb <= "101111";
					when "101000100001101" => rgb <= "101111";
					when "101000100001110" => rgb <= "101111";
					when "101000100001111" => rgb <= "101111";
					when "101000100010000" => rgb <= "101111";
					when "101000100010001" => rgb <= "101111";
					when "101000100010010" => rgb <= "101111";
					when "101000100010011" => rgb <= "101111";
					when "101000100010100" => rgb <= "101111";
					when "101000100010101" => rgb <= "101111";
					when "101000100010110" => rgb <= "101111";
					when "101000100010111" => rgb <= "101111";
					when "101000100011000" => rgb <= "101111";
					when "101000100011001" => rgb <= "101111";
					when "101000100011010" => rgb <= "101111";
					when "101000100011011" => rgb <= "101111";
					when "101000100011100" => rgb <= "101111";
					when "101000100011101" => rgb <= "101111";
					when "101000100011110" => rgb <= "101111";
					when "101000100011111" => rgb <= "101111";
					when "101000100100000" => rgb <= "000000";
					when "101000100100001" => rgb <= "000000";
					when "101000100100010" => rgb <= "100100";
					when "101000100100011" => rgb <= "100100";
					when "101000100100100" => rgb <= "100100";
					when "101000100100101" => rgb <= "100100";
					when "101000100100110" => rgb <= "100100";
					when "101000100100111" => rgb <= "100100";
					when "101000100101000" => rgb <= "100100";
					when "101000100101001" => rgb <= "100100";
					when "101000100101010" => rgb <= "100100";
					when "101000100101011" => rgb <= "100100";
					when "101000100101100" => rgb <= "000000";
					when "101000100101101" => rgb <= "000000";
					when "101000100101110" => rgb <= "100100";
					when "101000100101111" => rgb <= "100100";
					when "101000100110000" => rgb <= "100100";
					when "101000100110001" => rgb <= "100100";
					when "101000100110010" => rgb <= "010000";
					when "101000100110011" => rgb <= "010000";
					when "101000100110100" => rgb <= "000000";
					when "101000100110101" => rgb <= "000000";
					when "101000100110110" => rgb <= "101111";
					when "101000100110111" => rgb <= "101111";
					when "101000100111000" => rgb <= "101111";
					when "101000100111001" => rgb <= "101111";
					when "101000100111010" => rgb <= "101111";
					when "101000100111011" => rgb <= "101111";
					when "101000100111100" => rgb <= "101111";
					when "101000100111101" => rgb <= "101111";
					when "101000100111110" => rgb <= "101111";
					when "101000100111111" => rgb <= "101111";
					when "101000101000000" => rgb <= "101111";
					when "101000101000001" => rgb <= "101111";
					when "101000101000010" => rgb <= "101111";
					when "101000101000011" => rgb <= "101111";
					when "101000101000100" => rgb <= "101111";
					when "101000101000101" => rgb <= "101111";
					when "101000101000110" => rgb <= "101111";
					when "101000101000111" => rgb <= "101111";
					when "101000101001000" => rgb <= "101111";
					when "101000101001001" => rgb <= "101111";
					when "101000101001010" => rgb <= "101111";
					when "101000101001011" => rgb <= "101111";
					when "101000101001100" => rgb <= "101111";
					when "101000101001101" => rgb <= "101111";
					when "101000101001110" => rgb <= "101111";
					when "101000101001111" => rgb <= "101111";
					when "101000101010000" => rgb <= "101111";
					when "101000101010001" => rgb <= "101111";
					when "101000101010010" => rgb <= "101111";
					when "101000101010011" => rgb <= "101111";
					when "101000101010100" => rgb <= "101111";
					when "101000101010101" => rgb <= "101111";
					when "101000101010110" => rgb <= "101111";
					when "101000101010111" => rgb <= "101111";
					when "101000101011000" => rgb <= "101111";
					when "101000101011001" => rgb <= "101111";
					when "101000101011010" => rgb <= "101111";
					when "101000101011011" => rgb <= "101111";
					when "101000101011100" => rgb <= "101111";
					when "101000101011101" => rgb <= "101111";
					when "101000101011110" => rgb <= "101111";
					when "101000101011111" => rgb <= "101111";
					when "101000101100000" => rgb <= "101111";
					when "101000101100001" => rgb <= "101111";
					when "101000101100010" => rgb <= "101111";
					when "101000101100011" => rgb <= "101111";
					when "101000101100100" => rgb <= "101111";
					when "101000101100101" => rgb <= "101111";
					when "101000101100110" => rgb <= "101111";
					when "101000101100111" => rgb <= "101111";
					when "101000101101000" => rgb <= "101111";
					when "101000101101001" => rgb <= "101111";
					when "101000101101010" => rgb <= "101111";
					when "101000101101011" => rgb <= "101111";
					when "101000101101100" => rgb <= "101111";
					when "101000101101101" => rgb <= "101111";
					when "101000101101110" => rgb <= "101111";
					when "101000101101111" => rgb <= "101111";
					when "101000101110000" => rgb <= "101111";
					when "101000101110001" => rgb <= "101111";
					when "101000101110010" => rgb <= "101111";
					when "101000101110011" => rgb <= "101111";
					when "101000101110100" => rgb <= "101111";
					when "101000101110101" => rgb <= "101111";
					when "101000101110110" => rgb <= "101111";
					when "101000101110111" => rgb <= "101111";
					when "101000101111000" => rgb <= "101111";
					when "101000101111001" => rgb <= "101111";
					when "101000101111010" => rgb <= "101111";
					when "101000101111011" => rgb <= "101111";
					when "101000101111100" => rgb <= "101111";
					when "101000101111101" => rgb <= "101111";
					when "101000101111110" => rgb <= "101111";
					when "101000101111111" => rgb <= "101111";
					when "101000110000000" => rgb <= "101111";
					when "101000110000001" => rgb <= "101111";
					when "101000110000010" => rgb <= "101111";
					when "101000110000011" => rgb <= "101111";
					when "101000110000100" => rgb <= "101111";
					when "101000110000101" => rgb <= "101111";
					when "101000110000110" => rgb <= "101111";
					when "101000110000111" => rgb <= "101111";
					when "101000110001000" => rgb <= "101111";
					when "101000110001001" => rgb <= "101111";
					when "101000110001010" => rgb <= "101111";
					when "101000110001011" => rgb <= "101111";
					when "101000110001100" => rgb <= "101111";
					when "101000110001101" => rgb <= "101111";
					when "101000110001110" => rgb <= "101111";
					when "101000110001111" => rgb <= "101111";
					when "101000110010000" => rgb <= "101111";
					when "101000110010001" => rgb <= "101111";
					when "101000110010010" => rgb <= "101111";
					when "101000110010011" => rgb <= "101111";
					when "101000110010100" => rgb <= "101111";
					when "101000110010101" => rgb <= "101111";
					when "101000110010110" => rgb <= "101111";
					when "101000110010111" => rgb <= "101111";
					when "101000110011000" => rgb <= "101111";
					when "101000110011001" => rgb <= "101111";
					when "101000110011010" => rgb <= "101111";
					when "101000110011011" => rgb <= "101111";
					when "101000110011100" => rgb <= "101111";
					when "101000110011101" => rgb <= "101111";
					when "101000110011110" => rgb <= "101111";
					when "101000110011111" => rgb <= "101111";
					when "101001000000000" => rgb <= "101111";
					when "101001000000001" => rgb <= "101111";
					when "101001000000010" => rgb <= "101111";
					when "101001000000011" => rgb <= "101111";
					when "101001000000100" => rgb <= "101111";
					when "101001000000101" => rgb <= "101111";
					when "101001000000110" => rgb <= "101111";
					when "101001000000111" => rgb <= "101111";
					when "101001000001000" => rgb <= "101111";
					when "101001000001001" => rgb <= "101111";
					when "101001000001010" => rgb <= "101111";
					when "101001000001011" => rgb <= "101111";
					when "101001000001100" => rgb <= "101111";
					when "101001000001101" => rgb <= "101111";
					when "101001000001110" => rgb <= "101111";
					when "101001000001111" => rgb <= "101111";
					when "101001000010000" => rgb <= "101111";
					when "101001000010001" => rgb <= "101111";
					when "101001000010010" => rgb <= "101111";
					when "101001000010011" => rgb <= "101111";
					when "101001000010100" => rgb <= "101111";
					when "101001000010101" => rgb <= "101111";
					when "101001000010110" => rgb <= "101111";
					when "101001000010111" => rgb <= "101111";
					when "101001000011000" => rgb <= "101111";
					when "101001000011001" => rgb <= "101111";
					when "101001000011010" => rgb <= "101111";
					when "101001000011011" => rgb <= "101111";
					when "101001000011100" => rgb <= "101111";
					when "101001000011101" => rgb <= "101111";
					when "101001000011110" => rgb <= "101111";
					when "101001000011111" => rgb <= "101111";
					when "101001000100000" => rgb <= "000000";
					when "101001000100001" => rgb <= "000000";
					when "101001000100010" => rgb <= "100100";
					when "101001000100011" => rgb <= "100100";
					when "101001000100100" => rgb <= "100100";
					when "101001000100101" => rgb <= "100100";
					when "101001000100110" => rgb <= "100100";
					when "101001000100111" => rgb <= "100100";
					when "101001000101000" => rgb <= "100100";
					when "101001000101001" => rgb <= "100100";
					when "101001000101010" => rgb <= "000000";
					when "101001000101011" => rgb <= "000000";
					when "101001000101100" => rgb <= "000000";
					when "101001000101101" => rgb <= "000000";
					when "101001000101110" => rgb <= "000000";
					when "101001000101111" => rgb <= "000000";
					when "101001000110000" => rgb <= "100100";
					when "101001000110001" => rgb <= "100100";
					when "101001000110010" => rgb <= "010000";
					when "101001000110011" => rgb <= "010000";
					when "101001000110100" => rgb <= "000000";
					when "101001000110101" => rgb <= "000000";
					when "101001000110110" => rgb <= "101111";
					when "101001000110111" => rgb <= "101111";
					when "101001000111000" => rgb <= "101111";
					when "101001000111001" => rgb <= "101111";
					when "101001000111010" => rgb <= "101111";
					when "101001000111011" => rgb <= "101111";
					when "101001000111100" => rgb <= "101111";
					when "101001000111101" => rgb <= "101111";
					when "101001000111110" => rgb <= "101111";
					when "101001000111111" => rgb <= "101111";
					when "101001001000000" => rgb <= "101111";
					when "101001001000001" => rgb <= "101111";
					when "101001001000010" => rgb <= "101111";
					when "101001001000011" => rgb <= "101111";
					when "101001001000100" => rgb <= "101111";
					when "101001001000101" => rgb <= "101111";
					when "101001001000110" => rgb <= "101111";
					when "101001001000111" => rgb <= "101111";
					when "101001001001000" => rgb <= "101111";
					when "101001001001001" => rgb <= "101111";
					when "101001001001010" => rgb <= "101111";
					when "101001001001011" => rgb <= "101111";
					when "101001001001100" => rgb <= "101111";
					when "101001001001101" => rgb <= "101111";
					when "101001001001110" => rgb <= "101111";
					when "101001001001111" => rgb <= "101111";
					when "101001001010000" => rgb <= "101111";
					when "101001001010001" => rgb <= "101111";
					when "101001001010010" => rgb <= "101111";
					when "101001001010011" => rgb <= "101111";
					when "101001001010100" => rgb <= "101111";
					when "101001001010101" => rgb <= "101111";
					when "101001001010110" => rgb <= "101111";
					when "101001001010111" => rgb <= "101111";
					when "101001001011000" => rgb <= "101111";
					when "101001001011001" => rgb <= "101111";
					when "101001001011010" => rgb <= "101111";
					when "101001001011011" => rgb <= "101111";
					when "101001001011100" => rgb <= "101111";
					when "101001001011101" => rgb <= "101111";
					when "101001001011110" => rgb <= "101111";
					when "101001001011111" => rgb <= "101111";
					when "101001001100000" => rgb <= "101111";
					when "101001001100001" => rgb <= "101111";
					when "101001001100010" => rgb <= "101111";
					when "101001001100011" => rgb <= "101111";
					when "101001001100100" => rgb <= "101111";
					when "101001001100101" => rgb <= "101111";
					when "101001001100110" => rgb <= "101111";
					when "101001001100111" => rgb <= "101111";
					when "101001001101000" => rgb <= "101111";
					when "101001001101001" => rgb <= "101111";
					when "101001001101010" => rgb <= "101111";
					when "101001001101011" => rgb <= "101111";
					when "101001001101100" => rgb <= "101111";
					when "101001001101101" => rgb <= "101111";
					when "101001001101110" => rgb <= "101111";
					when "101001001101111" => rgb <= "101111";
					when "101001001110000" => rgb <= "101111";
					when "101001001110001" => rgb <= "101111";
					when "101001001110010" => rgb <= "101111";
					when "101001001110011" => rgb <= "101111";
					when "101001001110100" => rgb <= "101111";
					when "101001001110101" => rgb <= "101111";
					when "101001001110110" => rgb <= "101111";
					when "101001001110111" => rgb <= "101111";
					when "101001001111000" => rgb <= "101111";
					when "101001001111001" => rgb <= "101111";
					when "101001001111010" => rgb <= "101111";
					when "101001001111011" => rgb <= "101111";
					when "101001001111100" => rgb <= "101111";
					when "101001001111101" => rgb <= "101111";
					when "101001001111110" => rgb <= "101111";
					when "101001001111111" => rgb <= "101111";
					when "101001010000000" => rgb <= "101111";
					when "101001010000001" => rgb <= "101111";
					when "101001010000010" => rgb <= "101111";
					when "101001010000011" => rgb <= "101111";
					when "101001010000100" => rgb <= "101111";
					when "101001010000101" => rgb <= "101111";
					when "101001010000110" => rgb <= "101111";
					when "101001010000111" => rgb <= "101111";
					when "101001010001000" => rgb <= "101111";
					when "101001010001001" => rgb <= "101111";
					when "101001010001010" => rgb <= "101111";
					when "101001010001011" => rgb <= "101111";
					when "101001010001100" => rgb <= "101111";
					when "101001010001101" => rgb <= "101111";
					when "101001010001110" => rgb <= "101111";
					when "101001010001111" => rgb <= "101111";
					when "101001010010000" => rgb <= "101111";
					when "101001010010001" => rgb <= "101111";
					when "101001010010010" => rgb <= "101111";
					when "101001010010011" => rgb <= "101111";
					when "101001010010100" => rgb <= "101111";
					when "101001010010101" => rgb <= "101111";
					when "101001010010110" => rgb <= "101111";
					when "101001010010111" => rgb <= "101111";
					when "101001010011000" => rgb <= "101111";
					when "101001010011001" => rgb <= "101111";
					when "101001010011010" => rgb <= "101111";
					when "101001010011011" => rgb <= "101111";
					when "101001010011100" => rgb <= "101111";
					when "101001010011101" => rgb <= "101111";
					when "101001010011110" => rgb <= "101111";
					when "101001010011111" => rgb <= "101111";
					when "101001100000000" => rgb <= "101111";
					when "101001100000001" => rgb <= "101111";
					when "101001100000010" => rgb <= "101111";
					when "101001100000011" => rgb <= "101111";
					when "101001100000100" => rgb <= "101111";
					when "101001100000101" => rgb <= "101111";
					when "101001100000110" => rgb <= "101111";
					when "101001100000111" => rgb <= "101111";
					when "101001100001000" => rgb <= "101111";
					when "101001100001001" => rgb <= "101111";
					when "101001100001010" => rgb <= "101111";
					when "101001100001011" => rgb <= "101111";
					when "101001100001100" => rgb <= "101111";
					when "101001100001101" => rgb <= "101111";
					when "101001100001110" => rgb <= "101111";
					when "101001100001111" => rgb <= "101111";
					when "101001100010000" => rgb <= "101111";
					when "101001100010001" => rgb <= "101111";
					when "101001100010010" => rgb <= "101111";
					when "101001100010011" => rgb <= "101111";
					when "101001100010100" => rgb <= "101111";
					when "101001100010101" => rgb <= "101111";
					when "101001100010110" => rgb <= "101111";
					when "101001100010111" => rgb <= "101111";
					when "101001100011000" => rgb <= "101111";
					when "101001100011001" => rgb <= "101111";
					when "101001100011010" => rgb <= "101111";
					when "101001100011011" => rgb <= "101111";
					when "101001100011100" => rgb <= "101111";
					when "101001100011101" => rgb <= "101111";
					when "101001100011110" => rgb <= "101111";
					when "101001100011111" => rgb <= "101111";
					when "101001100100000" => rgb <= "000000";
					when "101001100100001" => rgb <= "000000";
					when "101001100100010" => rgb <= "100100";
					when "101001100100011" => rgb <= "100100";
					when "101001100100100" => rgb <= "100100";
					when "101001100100101" => rgb <= "100100";
					when "101001100100110" => rgb <= "100100";
					when "101001100100111" => rgb <= "100100";
					when "101001100101000" => rgb <= "100100";
					when "101001100101001" => rgb <= "100100";
					when "101001100101010" => rgb <= "000000";
					when "101001100101011" => rgb <= "000000";
					when "101001100101100" => rgb <= "000000";
					when "101001100101101" => rgb <= "000000";
					when "101001100101110" => rgb <= "000000";
					when "101001100101111" => rgb <= "000000";
					when "101001100110000" => rgb <= "100100";
					when "101001100110001" => rgb <= "100100";
					when "101001100110010" => rgb <= "010000";
					when "101001100110011" => rgb <= "010000";
					when "101001100110100" => rgb <= "000000";
					when "101001100110101" => rgb <= "000000";
					when "101001100110110" => rgb <= "101111";
					when "101001100110111" => rgb <= "101111";
					when "101001100111000" => rgb <= "101111";
					when "101001100111001" => rgb <= "101111";
					when "101001100111010" => rgb <= "101111";
					when "101001100111011" => rgb <= "101111";
					when "101001100111100" => rgb <= "101111";
					when "101001100111101" => rgb <= "101111";
					when "101001100111110" => rgb <= "101111";
					when "101001100111111" => rgb <= "101111";
					when "101001101000000" => rgb <= "101111";
					when "101001101000001" => rgb <= "101111";
					when "101001101000010" => rgb <= "101111";
					when "101001101000011" => rgb <= "101111";
					when "101001101000100" => rgb <= "101111";
					when "101001101000101" => rgb <= "101111";
					when "101001101000110" => rgb <= "101111";
					when "101001101000111" => rgb <= "101111";
					when "101001101001000" => rgb <= "101111";
					when "101001101001001" => rgb <= "101111";
					when "101001101001010" => rgb <= "101111";
					when "101001101001011" => rgb <= "101111";
					when "101001101001100" => rgb <= "101111";
					when "101001101001101" => rgb <= "101111";
					when "101001101001110" => rgb <= "101111";
					when "101001101001111" => rgb <= "101111";
					when "101001101010000" => rgb <= "101111";
					when "101001101010001" => rgb <= "101111";
					when "101001101010010" => rgb <= "101111";
					when "101001101010011" => rgb <= "101111";
					when "101001101010100" => rgb <= "101111";
					when "101001101010101" => rgb <= "101111";
					when "101001101010110" => rgb <= "101111";
					when "101001101010111" => rgb <= "101111";
					when "101001101011000" => rgb <= "101111";
					when "101001101011001" => rgb <= "101111";
					when "101001101011010" => rgb <= "101111";
					when "101001101011011" => rgb <= "101111";
					when "101001101011100" => rgb <= "101111";
					when "101001101011101" => rgb <= "101111";
					when "101001101011110" => rgb <= "101111";
					when "101001101011111" => rgb <= "101111";
					when "101001101100000" => rgb <= "101111";
					when "101001101100001" => rgb <= "101111";
					when "101001101100010" => rgb <= "101111";
					when "101001101100011" => rgb <= "101111";
					when "101001101100100" => rgb <= "101111";
					when "101001101100101" => rgb <= "101111";
					when "101001101100110" => rgb <= "101111";
					when "101001101100111" => rgb <= "101111";
					when "101001101101000" => rgb <= "101111";
					when "101001101101001" => rgb <= "101111";
					when "101001101101010" => rgb <= "101111";
					when "101001101101011" => rgb <= "101111";
					when "101001101101100" => rgb <= "101111";
					when "101001101101101" => rgb <= "101111";
					when "101001101101110" => rgb <= "101111";
					when "101001101101111" => rgb <= "101111";
					when "101001101110000" => rgb <= "101111";
					when "101001101110001" => rgb <= "101111";
					when "101001101110010" => rgb <= "101111";
					when "101001101110011" => rgb <= "101111";
					when "101001101110100" => rgb <= "101111";
					when "101001101110101" => rgb <= "101111";
					when "101001101110110" => rgb <= "101111";
					when "101001101110111" => rgb <= "101111";
					when "101001101111000" => rgb <= "101111";
					when "101001101111001" => rgb <= "101111";
					when "101001101111010" => rgb <= "101111";
					when "101001101111011" => rgb <= "101111";
					when "101001101111100" => rgb <= "101111";
					when "101001101111101" => rgb <= "101111";
					when "101001101111110" => rgb <= "101111";
					when "101001101111111" => rgb <= "101111";
					when "101001110000000" => rgb <= "101111";
					when "101001110000001" => rgb <= "101111";
					when "101001110000010" => rgb <= "101111";
					when "101001110000011" => rgb <= "101111";
					when "101001110000100" => rgb <= "101111";
					when "101001110000101" => rgb <= "101111";
					when "101001110000110" => rgb <= "101111";
					when "101001110000111" => rgb <= "101111";
					when "101001110001000" => rgb <= "101111";
					when "101001110001001" => rgb <= "101111";
					when "101001110001010" => rgb <= "101111";
					when "101001110001011" => rgb <= "101111";
					when "101001110001100" => rgb <= "101111";
					when "101001110001101" => rgb <= "101111";
					when "101001110001110" => rgb <= "101111";
					when "101001110001111" => rgb <= "101111";
					when "101001110010000" => rgb <= "101111";
					when "101001110010001" => rgb <= "101111";
					when "101001110010010" => rgb <= "101111";
					when "101001110010011" => rgb <= "101111";
					when "101001110010100" => rgb <= "101111";
					when "101001110010101" => rgb <= "101111";
					when "101001110010110" => rgb <= "101111";
					when "101001110010111" => rgb <= "101111";
					when "101001110011000" => rgb <= "101111";
					when "101001110011001" => rgb <= "101111";
					when "101001110011010" => rgb <= "101111";
					when "101001110011011" => rgb <= "101111";
					when "101001110011100" => rgb <= "101111";
					when "101001110011101" => rgb <= "101111";
					when "101001110011110" => rgb <= "101111";
					when "101001110011111" => rgb <= "101111";
					when "101010000000000" => rgb <= "101111";
					when "101010000000001" => rgb <= "101111";
					when "101010000000010" => rgb <= "101111";
					when "101010000000011" => rgb <= "101111";
					when "101010000000100" => rgb <= "101111";
					when "101010000000101" => rgb <= "101111";
					when "101010000000110" => rgb <= "101111";
					when "101010000000111" => rgb <= "101111";
					when "101010000001000" => rgb <= "101111";
					when "101010000001001" => rgb <= "101111";
					when "101010000001010" => rgb <= "101111";
					when "101010000001011" => rgb <= "101111";
					when "101010000001100" => rgb <= "101111";
					when "101010000001101" => rgb <= "101111";
					when "101010000001110" => rgb <= "101111";
					when "101010000001111" => rgb <= "101111";
					when "101010000010000" => rgb <= "101111";
					when "101010000010001" => rgb <= "101111";
					when "101010000010010" => rgb <= "101111";
					when "101010000010011" => rgb <= "101111";
					when "101010000010100" => rgb <= "101111";
					when "101010000010101" => rgb <= "101111";
					when "101010000010110" => rgb <= "101111";
					when "101010000010111" => rgb <= "101111";
					when "101010000011000" => rgb <= "101111";
					when "101010000011001" => rgb <= "101111";
					when "101010000011010" => rgb <= "101111";
					when "101010000011011" => rgb <= "101111";
					when "101010000011100" => rgb <= "101111";
					when "101010000011101" => rgb <= "101111";
					when "101010000011110" => rgb <= "101111";
					when "101010000011111" => rgb <= "101111";
					when "101010000100000" => rgb <= "000000";
					when "101010000100001" => rgb <= "000000";
					when "101010000100010" => rgb <= "100100";
					when "101010000100011" => rgb <= "100100";
					when "101010000100100" => rgb <= "100100";
					when "101010000100101" => rgb <= "100100";
					when "101010000100110" => rgb <= "100100";
					when "101010000100111" => rgb <= "100100";
					when "101010000101000" => rgb <= "100100";
					when "101010000101001" => rgb <= "100100";
					when "101010000101010" => rgb <= "100100";
					when "101010000101011" => rgb <= "100100";
					when "101010000101100" => rgb <= "000000";
					when "101010000101101" => rgb <= "000000";
					when "101010000101110" => rgb <= "100100";
					when "101010000101111" => rgb <= "100100";
					when "101010000110000" => rgb <= "100100";
					when "101010000110001" => rgb <= "100100";
					when "101010000110010" => rgb <= "010000";
					when "101010000110011" => rgb <= "010000";
					when "101010000110100" => rgb <= "000000";
					when "101010000110101" => rgb <= "000000";
					when "101010000110110" => rgb <= "101111";
					when "101010000110111" => rgb <= "101111";
					when "101010000111000" => rgb <= "101111";
					when "101010000111001" => rgb <= "101111";
					when "101010000111010" => rgb <= "101111";
					when "101010000111011" => rgb <= "101111";
					when "101010000111100" => rgb <= "101111";
					when "101010000111101" => rgb <= "101111";
					when "101010000111110" => rgb <= "101111";
					when "101010000111111" => rgb <= "101111";
					when "101010001000000" => rgb <= "101111";
					when "101010001000001" => rgb <= "101111";
					when "101010001000010" => rgb <= "101111";
					when "101010001000011" => rgb <= "101111";
					when "101010001000100" => rgb <= "101111";
					when "101010001000101" => rgb <= "101111";
					when "101010001000110" => rgb <= "101111";
					when "101010001000111" => rgb <= "101111";
					when "101010001001000" => rgb <= "101111";
					when "101010001001001" => rgb <= "101111";
					when "101010001001010" => rgb <= "101111";
					when "101010001001011" => rgb <= "101111";
					when "101010001001100" => rgb <= "101111";
					when "101010001001101" => rgb <= "101111";
					when "101010001001110" => rgb <= "101111";
					when "101010001001111" => rgb <= "101111";
					when "101010001010000" => rgb <= "101111";
					when "101010001010001" => rgb <= "101111";
					when "101010001010010" => rgb <= "101111";
					when "101010001010011" => rgb <= "101111";
					when "101010001010100" => rgb <= "101111";
					when "101010001010101" => rgb <= "101111";
					when "101010001010110" => rgb <= "101111";
					when "101010001010111" => rgb <= "101111";
					when "101010001011000" => rgb <= "101111";
					when "101010001011001" => rgb <= "101111";
					when "101010001011010" => rgb <= "101111";
					when "101010001011011" => rgb <= "101111";
					when "101010001011100" => rgb <= "101111";
					when "101010001011101" => rgb <= "101111";
					when "101010001011110" => rgb <= "101111";
					when "101010001011111" => rgb <= "101111";
					when "101010001100000" => rgb <= "101111";
					when "101010001100001" => rgb <= "101111";
					when "101010001100010" => rgb <= "101111";
					when "101010001100011" => rgb <= "101111";
					when "101010001100100" => rgb <= "101111";
					when "101010001100101" => rgb <= "101111";
					when "101010001100110" => rgb <= "101111";
					when "101010001100111" => rgb <= "101111";
					when "101010001101000" => rgb <= "101111";
					when "101010001101001" => rgb <= "101111";
					when "101010001101010" => rgb <= "101111";
					when "101010001101011" => rgb <= "101111";
					when "101010001101100" => rgb <= "101111";
					when "101010001101101" => rgb <= "101111";
					when "101010001101110" => rgb <= "101111";
					when "101010001101111" => rgb <= "101111";
					when "101010001110000" => rgb <= "101111";
					when "101010001110001" => rgb <= "101111";
					when "101010001110010" => rgb <= "101111";
					when "101010001110011" => rgb <= "101111";
					when "101010001110100" => rgb <= "101111";
					when "101010001110101" => rgb <= "101111";
					when "101010001110110" => rgb <= "101111";
					when "101010001110111" => rgb <= "101111";
					when "101010001111000" => rgb <= "101111";
					when "101010001111001" => rgb <= "101111";
					when "101010001111010" => rgb <= "101111";
					when "101010001111011" => rgb <= "101111";
					when "101010001111100" => rgb <= "101111";
					when "101010001111101" => rgb <= "101111";
					when "101010001111110" => rgb <= "101111";
					when "101010001111111" => rgb <= "101111";
					when "101010010000000" => rgb <= "101111";
					when "101010010000001" => rgb <= "101111";
					when "101010010000010" => rgb <= "101111";
					when "101010010000011" => rgb <= "101111";
					when "101010010000100" => rgb <= "101111";
					when "101010010000101" => rgb <= "101111";
					when "101010010000110" => rgb <= "101111";
					when "101010010000111" => rgb <= "101111";
					when "101010010001000" => rgb <= "101111";
					when "101010010001001" => rgb <= "101111";
					when "101010010001010" => rgb <= "101111";
					when "101010010001011" => rgb <= "101111";
					when "101010010001100" => rgb <= "101111";
					when "101010010001101" => rgb <= "101111";
					when "101010010001110" => rgb <= "101111";
					when "101010010001111" => rgb <= "101111";
					when "101010010010000" => rgb <= "101111";
					when "101010010010001" => rgb <= "101111";
					when "101010010010010" => rgb <= "101111";
					when "101010010010011" => rgb <= "101111";
					when "101010010010100" => rgb <= "101111";
					when "101010010010101" => rgb <= "101111";
					when "101010010010110" => rgb <= "101111";
					when "101010010010111" => rgb <= "101111";
					when "101010010011000" => rgb <= "101111";
					when "101010010011001" => rgb <= "101111";
					when "101010010011010" => rgb <= "101111";
					when "101010010011011" => rgb <= "101111";
					when "101010010011100" => rgb <= "101111";
					when "101010010011101" => rgb <= "101111";
					when "101010010011110" => rgb <= "101111";
					when "101010010011111" => rgb <= "101111";
					when "101010100000000" => rgb <= "101111";
					when "101010100000001" => rgb <= "101111";
					when "101010100000010" => rgb <= "101111";
					when "101010100000011" => rgb <= "101111";
					when "101010100000100" => rgb <= "101111";
					when "101010100000101" => rgb <= "101111";
					when "101010100000110" => rgb <= "101111";
					when "101010100000111" => rgb <= "101111";
					when "101010100001000" => rgb <= "101111";
					when "101010100001001" => rgb <= "101111";
					when "101010100001010" => rgb <= "101111";
					when "101010100001011" => rgb <= "101111";
					when "101010100001100" => rgb <= "101111";
					when "101010100001101" => rgb <= "101111";
					when "101010100001110" => rgb <= "101111";
					when "101010100001111" => rgb <= "101111";
					when "101010100010000" => rgb <= "101111";
					when "101010100010001" => rgb <= "101111";
					when "101010100010010" => rgb <= "101111";
					when "101010100010011" => rgb <= "101111";
					when "101010100010100" => rgb <= "101111";
					when "101010100010101" => rgb <= "101111";
					when "101010100010110" => rgb <= "101111";
					when "101010100010111" => rgb <= "101111";
					when "101010100011000" => rgb <= "101111";
					when "101010100011001" => rgb <= "101111";
					when "101010100011010" => rgb <= "101111";
					when "101010100011011" => rgb <= "101111";
					when "101010100011100" => rgb <= "101111";
					when "101010100011101" => rgb <= "101111";
					when "101010100011110" => rgb <= "101111";
					when "101010100011111" => rgb <= "101111";
					when "101010100100000" => rgb <= "000000";
					when "101010100100001" => rgb <= "000000";
					when "101010100100010" => rgb <= "100100";
					when "101010100100011" => rgb <= "100100";
					when "101010100100100" => rgb <= "100100";
					when "101010100100101" => rgb <= "100100";
					when "101010100100110" => rgb <= "100100";
					when "101010100100111" => rgb <= "100100";
					when "101010100101000" => rgb <= "100100";
					when "101010100101001" => rgb <= "100100";
					when "101010100101010" => rgb <= "100100";
					when "101010100101011" => rgb <= "100100";
					when "101010100101100" => rgb <= "000000";
					when "101010100101101" => rgb <= "000000";
					when "101010100101110" => rgb <= "100100";
					when "101010100101111" => rgb <= "100100";
					when "101010100110000" => rgb <= "100100";
					when "101010100110001" => rgb <= "100100";
					when "101010100110010" => rgb <= "010000";
					when "101010100110011" => rgb <= "010000";
					when "101010100110100" => rgb <= "000000";
					when "101010100110101" => rgb <= "000000";
					when "101010100110110" => rgb <= "101111";
					when "101010100110111" => rgb <= "101111";
					when "101010100111000" => rgb <= "101111";
					when "101010100111001" => rgb <= "101111";
					when "101010100111010" => rgb <= "101111";
					when "101010100111011" => rgb <= "101111";
					when "101010100111100" => rgb <= "101111";
					when "101010100111101" => rgb <= "101111";
					when "101010100111110" => rgb <= "101111";
					when "101010100111111" => rgb <= "101111";
					when "101010101000000" => rgb <= "101111";
					when "101010101000001" => rgb <= "101111";
					when "101010101000010" => rgb <= "101111";
					when "101010101000011" => rgb <= "101111";
					when "101010101000100" => rgb <= "101111";
					when "101010101000101" => rgb <= "101111";
					when "101010101000110" => rgb <= "101111";
					when "101010101000111" => rgb <= "101111";
					when "101010101001000" => rgb <= "101111";
					when "101010101001001" => rgb <= "101111";
					when "101010101001010" => rgb <= "101111";
					when "101010101001011" => rgb <= "101111";
					when "101010101001100" => rgb <= "101111";
					when "101010101001101" => rgb <= "101111";
					when "101010101001110" => rgb <= "101111";
					when "101010101001111" => rgb <= "101111";
					when "101010101010000" => rgb <= "101111";
					when "101010101010001" => rgb <= "101111";
					when "101010101010010" => rgb <= "101111";
					when "101010101010011" => rgb <= "101111";
					when "101010101010100" => rgb <= "101111";
					when "101010101010101" => rgb <= "101111";
					when "101010101010110" => rgb <= "101111";
					when "101010101010111" => rgb <= "101111";
					when "101010101011000" => rgb <= "101111";
					when "101010101011001" => rgb <= "101111";
					when "101010101011010" => rgb <= "101111";
					when "101010101011011" => rgb <= "101111";
					when "101010101011100" => rgb <= "101111";
					when "101010101011101" => rgb <= "101111";
					when "101010101011110" => rgb <= "101111";
					when "101010101011111" => rgb <= "101111";
					when "101010101100000" => rgb <= "101111";
					when "101010101100001" => rgb <= "101111";
					when "101010101100010" => rgb <= "101111";
					when "101010101100011" => rgb <= "101111";
					when "101010101100100" => rgb <= "101111";
					when "101010101100101" => rgb <= "101111";
					when "101010101100110" => rgb <= "101111";
					when "101010101100111" => rgb <= "101111";
					when "101010101101000" => rgb <= "101111";
					when "101010101101001" => rgb <= "101111";
					when "101010101101010" => rgb <= "101111";
					when "101010101101011" => rgb <= "101111";
					when "101010101101100" => rgb <= "101111";
					when "101010101101101" => rgb <= "101111";
					when "101010101101110" => rgb <= "101111";
					when "101010101101111" => rgb <= "101111";
					when "101010101110000" => rgb <= "101111";
					when "101010101110001" => rgb <= "101111";
					when "101010101110010" => rgb <= "101111";
					when "101010101110011" => rgb <= "101111";
					when "101010101110100" => rgb <= "101111";
					when "101010101110101" => rgb <= "101111";
					when "101010101110110" => rgb <= "101111";
					when "101010101110111" => rgb <= "101111";
					when "101010101111000" => rgb <= "101111";
					when "101010101111001" => rgb <= "101111";
					when "101010101111010" => rgb <= "101111";
					when "101010101111011" => rgb <= "101111";
					when "101010101111100" => rgb <= "101111";
					when "101010101111101" => rgb <= "101111";
					when "101010101111110" => rgb <= "101111";
					when "101010101111111" => rgb <= "101111";
					when "101010110000000" => rgb <= "101111";
					when "101010110000001" => rgb <= "101111";
					when "101010110000010" => rgb <= "101111";
					when "101010110000011" => rgb <= "101111";
					when "101010110000100" => rgb <= "101111";
					when "101010110000101" => rgb <= "101111";
					when "101010110000110" => rgb <= "101111";
					when "101010110000111" => rgb <= "101111";
					when "101010110001000" => rgb <= "101111";
					when "101010110001001" => rgb <= "101111";
					when "101010110001010" => rgb <= "101111";
					when "101010110001011" => rgb <= "101111";
					when "101010110001100" => rgb <= "101111";
					when "101010110001101" => rgb <= "101111";
					when "101010110001110" => rgb <= "101111";
					when "101010110001111" => rgb <= "101111";
					when "101010110010000" => rgb <= "101111";
					when "101010110010001" => rgb <= "101111";
					when "101010110010010" => rgb <= "101111";
					when "101010110010011" => rgb <= "101111";
					when "101010110010100" => rgb <= "101111";
					when "101010110010101" => rgb <= "101111";
					when "101010110010110" => rgb <= "101111";
					when "101010110010111" => rgb <= "101111";
					when "101010110011000" => rgb <= "101111";
					when "101010110011001" => rgb <= "101111";
					when "101010110011010" => rgb <= "101111";
					when "101010110011011" => rgb <= "101111";
					when "101010110011100" => rgb <= "101111";
					when "101010110011101" => rgb <= "101111";
					when "101010110011110" => rgb <= "101111";
					when "101010110011111" => rgb <= "101111";
					when "101011000000000" => rgb <= "101111";
					when "101011000000001" => rgb <= "101111";
					when "101011000000010" => rgb <= "101111";
					when "101011000000011" => rgb <= "101111";
					when "101011000000100" => rgb <= "101111";
					when "101011000000101" => rgb <= "101111";
					when "101011000000110" => rgb <= "101111";
					when "101011000000111" => rgb <= "101111";
					when "101011000001000" => rgb <= "101111";
					when "101011000001001" => rgb <= "101111";
					when "101011000001010" => rgb <= "101111";
					when "101011000001011" => rgb <= "101111";
					when "101011000001100" => rgb <= "101111";
					when "101011000001101" => rgb <= "101111";
					when "101011000001110" => rgb <= "101111";
					when "101011000001111" => rgb <= "101111";
					when "101011000010000" => rgb <= "101111";
					when "101011000010001" => rgb <= "101111";
					when "101011000010010" => rgb <= "101111";
					when "101011000010011" => rgb <= "101111";
					when "101011000010100" => rgb <= "101111";
					when "101011000010101" => rgb <= "101111";
					when "101011000010110" => rgb <= "101111";
					when "101011000010111" => rgb <= "101111";
					when "101011000011000" => rgb <= "101111";
					when "101011000011001" => rgb <= "101111";
					when "101011000011010" => rgb <= "101111";
					when "101011000011011" => rgb <= "101111";
					when "101011000011100" => rgb <= "101111";
					when "101011000011101" => rgb <= "101111";
					when "101011000011110" => rgb <= "101111";
					when "101011000011111" => rgb <= "101111";
					when "101011000100000" => rgb <= "000000";
					when "101011000100001" => rgb <= "000000";
					when "101011000100010" => rgb <= "100100";
					when "101011000100011" => rgb <= "100100";
					when "101011000100100" => rgb <= "100100";
					when "101011000100101" => rgb <= "100100";
					when "101011000100110" => rgb <= "100100";
					when "101011000100111" => rgb <= "100100";
					when "101011000101000" => rgb <= "100100";
					when "101011000101001" => rgb <= "100100";
					when "101011000101010" => rgb <= "100100";
					when "101011000101011" => rgb <= "100100";
					when "101011000101100" => rgb <= "100100";
					when "101011000101101" => rgb <= "100100";
					when "101011000101110" => rgb <= "100100";
					when "101011000101111" => rgb <= "100100";
					when "101011000110000" => rgb <= "100100";
					when "101011000110001" => rgb <= "100100";
					when "101011000110010" => rgb <= "010000";
					when "101011000110011" => rgb <= "010000";
					when "101011000110100" => rgb <= "000000";
					when "101011000110101" => rgb <= "000000";
					when "101011000110110" => rgb <= "101111";
					when "101011000110111" => rgb <= "101111";
					when "101011000111000" => rgb <= "101111";
					when "101011000111001" => rgb <= "101111";
					when "101011000111010" => rgb <= "101111";
					when "101011000111011" => rgb <= "101111";
					when "101011000111100" => rgb <= "101111";
					when "101011000111101" => rgb <= "101111";
					when "101011000111110" => rgb <= "101111";
					when "101011000111111" => rgb <= "101111";
					when "101011001000000" => rgb <= "101111";
					when "101011001000001" => rgb <= "101111";
					when "101011001000010" => rgb <= "101111";
					when "101011001000011" => rgb <= "101111";
					when "101011001000100" => rgb <= "101111";
					when "101011001000101" => rgb <= "101111";
					when "101011001000110" => rgb <= "101111";
					when "101011001000111" => rgb <= "101111";
					when "101011001001000" => rgb <= "101111";
					when "101011001001001" => rgb <= "101111";
					when "101011001001010" => rgb <= "101111";
					when "101011001001011" => rgb <= "101111";
					when "101011001001100" => rgb <= "101111";
					when "101011001001101" => rgb <= "101111";
					when "101011001001110" => rgb <= "101111";
					when "101011001001111" => rgb <= "101111";
					when "101011001010000" => rgb <= "101111";
					when "101011001010001" => rgb <= "101111";
					when "101011001010010" => rgb <= "101111";
					when "101011001010011" => rgb <= "101111";
					when "101011001010100" => rgb <= "101111";
					when "101011001010101" => rgb <= "101111";
					when "101011001010110" => rgb <= "101111";
					when "101011001010111" => rgb <= "101111";
					when "101011001011000" => rgb <= "101111";
					when "101011001011001" => rgb <= "101111";
					when "101011001011010" => rgb <= "101111";
					when "101011001011011" => rgb <= "101111";
					when "101011001011100" => rgb <= "101111";
					when "101011001011101" => rgb <= "101111";
					when "101011001011110" => rgb <= "101111";
					when "101011001011111" => rgb <= "101111";
					when "101011001100000" => rgb <= "101111";
					when "101011001100001" => rgb <= "101111";
					when "101011001100010" => rgb <= "101111";
					when "101011001100011" => rgb <= "101111";
					when "101011001100100" => rgb <= "101111";
					when "101011001100101" => rgb <= "101111";
					when "101011001100110" => rgb <= "101111";
					when "101011001100111" => rgb <= "101111";
					when "101011001101000" => rgb <= "101111";
					when "101011001101001" => rgb <= "101111";
					when "101011001101010" => rgb <= "101111";
					when "101011001101011" => rgb <= "101111";
					when "101011001101100" => rgb <= "101111";
					when "101011001101101" => rgb <= "101111";
					when "101011001101110" => rgb <= "101111";
					when "101011001101111" => rgb <= "101111";
					when "101011001110000" => rgb <= "101111";
					when "101011001110001" => rgb <= "101111";
					when "101011001110010" => rgb <= "101111";
					when "101011001110011" => rgb <= "101111";
					when "101011001110100" => rgb <= "101111";
					when "101011001110101" => rgb <= "101111";
					when "101011001110110" => rgb <= "101111";
					when "101011001110111" => rgb <= "101111";
					when "101011001111000" => rgb <= "101111";
					when "101011001111001" => rgb <= "101111";
					when "101011001111010" => rgb <= "101111";
					when "101011001111011" => rgb <= "101111";
					when "101011001111100" => rgb <= "101111";
					when "101011001111101" => rgb <= "101111";
					when "101011001111110" => rgb <= "101111";
					when "101011001111111" => rgb <= "101111";
					when "101011010000000" => rgb <= "101111";
					when "101011010000001" => rgb <= "101111";
					when "101011010000010" => rgb <= "101111";
					when "101011010000011" => rgb <= "101111";
					when "101011010000100" => rgb <= "101111";
					when "101011010000101" => rgb <= "101111";
					when "101011010000110" => rgb <= "101111";
					when "101011010000111" => rgb <= "101111";
					when "101011010001000" => rgb <= "101111";
					when "101011010001001" => rgb <= "101111";
					when "101011010001010" => rgb <= "101111";
					when "101011010001011" => rgb <= "101111";
					when "101011010001100" => rgb <= "101111";
					when "101011010001101" => rgb <= "101111";
					when "101011010001110" => rgb <= "101111";
					when "101011010001111" => rgb <= "101111";
					when "101011010010000" => rgb <= "101111";
					when "101011010010001" => rgb <= "101111";
					when "101011010010010" => rgb <= "101111";
					when "101011010010011" => rgb <= "101111";
					when "101011010010100" => rgb <= "101111";
					when "101011010010101" => rgb <= "101111";
					when "101011010010110" => rgb <= "101111";
					when "101011010010111" => rgb <= "101111";
					when "101011010011000" => rgb <= "101111";
					when "101011010011001" => rgb <= "101111";
					when "101011010011010" => rgb <= "101111";
					when "101011010011011" => rgb <= "101111";
					when "101011010011100" => rgb <= "101111";
					when "101011010011101" => rgb <= "101111";
					when "101011010011110" => rgb <= "101111";
					when "101011010011111" => rgb <= "101111";
					when "101011100000000" => rgb <= "101111";
					when "101011100000001" => rgb <= "101111";
					when "101011100000010" => rgb <= "101111";
					when "101011100000011" => rgb <= "101111";
					when "101011100000100" => rgb <= "101111";
					when "101011100000101" => rgb <= "101111";
					when "101011100000110" => rgb <= "101111";
					when "101011100000111" => rgb <= "101111";
					when "101011100001000" => rgb <= "101111";
					when "101011100001001" => rgb <= "101111";
					when "101011100001010" => rgb <= "101111";
					when "101011100001011" => rgb <= "101111";
					when "101011100001100" => rgb <= "101111";
					when "101011100001101" => rgb <= "101111";
					when "101011100001110" => rgb <= "101111";
					when "101011100001111" => rgb <= "101111";
					when "101011100010000" => rgb <= "101111";
					when "101011100010001" => rgb <= "101111";
					when "101011100010010" => rgb <= "101111";
					when "101011100010011" => rgb <= "101111";
					when "101011100010100" => rgb <= "101111";
					when "101011100010101" => rgb <= "101111";
					when "101011100010110" => rgb <= "101111";
					when "101011100010111" => rgb <= "101111";
					when "101011100011000" => rgb <= "101111";
					when "101011100011001" => rgb <= "101111";
					when "101011100011010" => rgb <= "101111";
					when "101011100011011" => rgb <= "101111";
					when "101011100011100" => rgb <= "101111";
					when "101011100011101" => rgb <= "101111";
					when "101011100011110" => rgb <= "101111";
					when "101011100011111" => rgb <= "101111";
					when "101011100100000" => rgb <= "000000";
					when "101011100100001" => rgb <= "000000";
					when "101011100100010" => rgb <= "100100";
					when "101011100100011" => rgb <= "100100";
					when "101011100100100" => rgb <= "100100";
					when "101011100100101" => rgb <= "100100";
					when "101011100100110" => rgb <= "100100";
					when "101011100100111" => rgb <= "100100";
					when "101011100101000" => rgb <= "100100";
					when "101011100101001" => rgb <= "100100";
					when "101011100101010" => rgb <= "100100";
					when "101011100101011" => rgb <= "100100";
					when "101011100101100" => rgb <= "100100";
					when "101011100101101" => rgb <= "100100";
					when "101011100101110" => rgb <= "100100";
					when "101011100101111" => rgb <= "100100";
					when "101011100110000" => rgb <= "100100";
					when "101011100110001" => rgb <= "100100";
					when "101011100110010" => rgb <= "010000";
					when "101011100110011" => rgb <= "010000";
					when "101011100110100" => rgb <= "000000";
					when "101011100110101" => rgb <= "000000";
					when "101011100110110" => rgb <= "101111";
					when "101011100110111" => rgb <= "101111";
					when "101011100111000" => rgb <= "101111";
					when "101011100111001" => rgb <= "101111";
					when "101011100111010" => rgb <= "101111";
					when "101011100111011" => rgb <= "101111";
					when "101011100111100" => rgb <= "101111";
					when "101011100111101" => rgb <= "101111";
					when "101011100111110" => rgb <= "101111";
					when "101011100111111" => rgb <= "101111";
					when "101011101000000" => rgb <= "101111";
					when "101011101000001" => rgb <= "101111";
					when "101011101000010" => rgb <= "101111";
					when "101011101000011" => rgb <= "101111";
					when "101011101000100" => rgb <= "101111";
					when "101011101000101" => rgb <= "101111";
					when "101011101000110" => rgb <= "101111";
					when "101011101000111" => rgb <= "101111";
					when "101011101001000" => rgb <= "101111";
					when "101011101001001" => rgb <= "101111";
					when "101011101001010" => rgb <= "101111";
					when "101011101001011" => rgb <= "101111";
					when "101011101001100" => rgb <= "101111";
					when "101011101001101" => rgb <= "101111";
					when "101011101001110" => rgb <= "101111";
					when "101011101001111" => rgb <= "101111";
					when "101011101010000" => rgb <= "101111";
					when "101011101010001" => rgb <= "101111";
					when "101011101010010" => rgb <= "101111";
					when "101011101010011" => rgb <= "101111";
					when "101011101010100" => rgb <= "101111";
					when "101011101010101" => rgb <= "101111";
					when "101011101010110" => rgb <= "101111";
					when "101011101010111" => rgb <= "101111";
					when "101011101011000" => rgb <= "101111";
					when "101011101011001" => rgb <= "101111";
					when "101011101011010" => rgb <= "101111";
					when "101011101011011" => rgb <= "101111";
					when "101011101011100" => rgb <= "101111";
					when "101011101011101" => rgb <= "101111";
					when "101011101011110" => rgb <= "101111";
					when "101011101011111" => rgb <= "101111";
					when "101011101100000" => rgb <= "101111";
					when "101011101100001" => rgb <= "101111";
					when "101011101100010" => rgb <= "101111";
					when "101011101100011" => rgb <= "101111";
					when "101011101100100" => rgb <= "101111";
					when "101011101100101" => rgb <= "101111";
					when "101011101100110" => rgb <= "101111";
					when "101011101100111" => rgb <= "101111";
					when "101011101101000" => rgb <= "101111";
					when "101011101101001" => rgb <= "101111";
					when "101011101101010" => rgb <= "101111";
					when "101011101101011" => rgb <= "101111";
					when "101011101101100" => rgb <= "101111";
					when "101011101101101" => rgb <= "101111";
					when "101011101101110" => rgb <= "101111";
					when "101011101101111" => rgb <= "101111";
					when "101011101110000" => rgb <= "101111";
					when "101011101110001" => rgb <= "101111";
					when "101011101110010" => rgb <= "101111";
					when "101011101110011" => rgb <= "101111";
					when "101011101110100" => rgb <= "101111";
					when "101011101110101" => rgb <= "101111";
					when "101011101110110" => rgb <= "101111";
					when "101011101110111" => rgb <= "101111";
					when "101011101111000" => rgb <= "101111";
					when "101011101111001" => rgb <= "101111";
					when "101011101111010" => rgb <= "101111";
					when "101011101111011" => rgb <= "101111";
					when "101011101111100" => rgb <= "101111";
					when "101011101111101" => rgb <= "101111";
					when "101011101111110" => rgb <= "101111";
					when "101011101111111" => rgb <= "101111";
					when "101011110000000" => rgb <= "101111";
					when "101011110000001" => rgb <= "101111";
					when "101011110000010" => rgb <= "101111";
					when "101011110000011" => rgb <= "101111";
					when "101011110000100" => rgb <= "101111";
					when "101011110000101" => rgb <= "101111";
					when "101011110000110" => rgb <= "101111";
					when "101011110000111" => rgb <= "101111";
					when "101011110001000" => rgb <= "101111";
					when "101011110001001" => rgb <= "101111";
					when "101011110001010" => rgb <= "101111";
					when "101011110001011" => rgb <= "101111";
					when "101011110001100" => rgb <= "101111";
					when "101011110001101" => rgb <= "101111";
					when "101011110001110" => rgb <= "101111";
					when "101011110001111" => rgb <= "101111";
					when "101011110010000" => rgb <= "101111";
					when "101011110010001" => rgb <= "101111";
					when "101011110010010" => rgb <= "101111";
					when "101011110010011" => rgb <= "101111";
					when "101011110010100" => rgb <= "101111";
					when "101011110010101" => rgb <= "101111";
					when "101011110010110" => rgb <= "101111";
					when "101011110010111" => rgb <= "101111";
					when "101011110011000" => rgb <= "101111";
					when "101011110011001" => rgb <= "101111";
					when "101011110011010" => rgb <= "101111";
					when "101011110011011" => rgb <= "101111";
					when "101011110011100" => rgb <= "101111";
					when "101011110011101" => rgb <= "101111";
					when "101011110011110" => rgb <= "101111";
					when "101011110011111" => rgb <= "101111";
					when "101100000000000" => rgb <= "101111";
					when "101100000000001" => rgb <= "101111";
					when "101100000000010" => rgb <= "101111";
					when "101100000000011" => rgb <= "101111";
					when "101100000000100" => rgb <= "101111";
					when "101100000000101" => rgb <= "101111";
					when "101100000000110" => rgb <= "101111";
					when "101100000000111" => rgb <= "101111";
					when "101100000001000" => rgb <= "101111";
					when "101100000001001" => rgb <= "101111";
					when "101100000001010" => rgb <= "101111";
					when "101100000001011" => rgb <= "101111";
					when "101100000001100" => rgb <= "101111";
					when "101100000001101" => rgb <= "101111";
					when "101100000001110" => rgb <= "101111";
					when "101100000001111" => rgb <= "101111";
					when "101100000010000" => rgb <= "101111";
					when "101100000010001" => rgb <= "101111";
					when "101100000010010" => rgb <= "101111";
					when "101100000010011" => rgb <= "101111";
					when "101100000010100" => rgb <= "101111";
					when "101100000010101" => rgb <= "101111";
					when "101100000010110" => rgb <= "101111";
					when "101100000010111" => rgb <= "101111";
					when "101100000011000" => rgb <= "101111";
					when "101100000011001" => rgb <= "101111";
					when "101100000011010" => rgb <= "101111";
					when "101100000011011" => rgb <= "101111";
					when "101100000011100" => rgb <= "101111";
					when "101100000011101" => rgb <= "101111";
					when "101100000011110" => rgb <= "101111";
					when "101100000011111" => rgb <= "101111";
					when "101100000100000" => rgb <= "000000";
					when "101100000100001" => rgb <= "000000";
					when "101100000100010" => rgb <= "100100";
					when "101100000100011" => rgb <= "100100";
					when "101100000100100" => rgb <= "100100";
					when "101100000100101" => rgb <= "100100";
					when "101100000100110" => rgb <= "100100";
					when "101100000100111" => rgb <= "100100";
					when "101100000101000" => rgb <= "100100";
					when "101100000101001" => rgb <= "100100";
					when "101100000101010" => rgb <= "100100";
					when "101100000101011" => rgb <= "100100";
					when "101100000101100" => rgb <= "100100";
					when "101100000101101" => rgb <= "100100";
					when "101100000101110" => rgb <= "100100";
					when "101100000101111" => rgb <= "100100";
					when "101100000110000" => rgb <= "100100";
					when "101100000110001" => rgb <= "100100";
					when "101100000110010" => rgb <= "010000";
					when "101100000110011" => rgb <= "010000";
					when "101100000110100" => rgb <= "000000";
					when "101100000110101" => rgb <= "000000";
					when "101100000110110" => rgb <= "101111";
					when "101100000110111" => rgb <= "101111";
					when "101100000111000" => rgb <= "101111";
					when "101100000111001" => rgb <= "101111";
					when "101100000111010" => rgb <= "101111";
					when "101100000111011" => rgb <= "101111";
					when "101100000111100" => rgb <= "101111";
					when "101100000111101" => rgb <= "101111";
					when "101100000111110" => rgb <= "101111";
					when "101100000111111" => rgb <= "101111";
					when "101100001000000" => rgb <= "101111";
					when "101100001000001" => rgb <= "101111";
					when "101100001000010" => rgb <= "101111";
					when "101100001000011" => rgb <= "101111";
					when "101100001000100" => rgb <= "101111";
					when "101100001000101" => rgb <= "101111";
					when "101100001000110" => rgb <= "101111";
					when "101100001000111" => rgb <= "101111";
					when "101100001001000" => rgb <= "101111";
					when "101100001001001" => rgb <= "101111";
					when "101100001001010" => rgb <= "101111";
					when "101100001001011" => rgb <= "101111";
					when "101100001001100" => rgb <= "101111";
					when "101100001001101" => rgb <= "101111";
					when "101100001001110" => rgb <= "101111";
					when "101100001001111" => rgb <= "101111";
					when "101100001010000" => rgb <= "101111";
					when "101100001010001" => rgb <= "101111";
					when "101100001010010" => rgb <= "101111";
					when "101100001010011" => rgb <= "101111";
					when "101100001010100" => rgb <= "101111";
					when "101100001010101" => rgb <= "101111";
					when "101100001010110" => rgb <= "101111";
					when "101100001010111" => rgb <= "101111";
					when "101100001011000" => rgb <= "101111";
					when "101100001011001" => rgb <= "101111";
					when "101100001011010" => rgb <= "101111";
					when "101100001011011" => rgb <= "101111";
					when "101100001011100" => rgb <= "101111";
					when "101100001011101" => rgb <= "101111";
					when "101100001011110" => rgb <= "101111";
					when "101100001011111" => rgb <= "101111";
					when "101100001100000" => rgb <= "101111";
					when "101100001100001" => rgb <= "101111";
					when "101100001100010" => rgb <= "101111";
					when "101100001100011" => rgb <= "101111";
					when "101100001100100" => rgb <= "101111";
					when "101100001100101" => rgb <= "101111";
					when "101100001100110" => rgb <= "101111";
					when "101100001100111" => rgb <= "101111";
					when "101100001101000" => rgb <= "101111";
					when "101100001101001" => rgb <= "101111";
					when "101100001101010" => rgb <= "101111";
					when "101100001101011" => rgb <= "101111";
					when "101100001101100" => rgb <= "101111";
					when "101100001101101" => rgb <= "101111";
					when "101100001101110" => rgb <= "101111";
					when "101100001101111" => rgb <= "101111";
					when "101100001110000" => rgb <= "101111";
					when "101100001110001" => rgb <= "101111";
					when "101100001110010" => rgb <= "101111";
					when "101100001110011" => rgb <= "101111";
					when "101100001110100" => rgb <= "101111";
					when "101100001110101" => rgb <= "101111";
					when "101100001110110" => rgb <= "101111";
					when "101100001110111" => rgb <= "101111";
					when "101100001111000" => rgb <= "101111";
					when "101100001111001" => rgb <= "101111";
					when "101100001111010" => rgb <= "101111";
					when "101100001111011" => rgb <= "101111";
					when "101100001111100" => rgb <= "101111";
					when "101100001111101" => rgb <= "101111";
					when "101100001111110" => rgb <= "101111";
					when "101100001111111" => rgb <= "101111";
					when "101100010000000" => rgb <= "101111";
					when "101100010000001" => rgb <= "101111";
					when "101100010000010" => rgb <= "101111";
					when "101100010000011" => rgb <= "101111";
					when "101100010000100" => rgb <= "101111";
					when "101100010000101" => rgb <= "101111";
					when "101100010000110" => rgb <= "101111";
					when "101100010000111" => rgb <= "101111";
					when "101100010001000" => rgb <= "101111";
					when "101100010001001" => rgb <= "101111";
					when "101100010001010" => rgb <= "101111";
					when "101100010001011" => rgb <= "101111";
					when "101100010001100" => rgb <= "101111";
					when "101100010001101" => rgb <= "101111";
					when "101100010001110" => rgb <= "101111";
					when "101100010001111" => rgb <= "101111";
					when "101100010010000" => rgb <= "101111";
					when "101100010010001" => rgb <= "101111";
					when "101100010010010" => rgb <= "101111";
					when "101100010010011" => rgb <= "101111";
					when "101100010010100" => rgb <= "101111";
					when "101100010010101" => rgb <= "101111";
					when "101100010010110" => rgb <= "101111";
					when "101100010010111" => rgb <= "101111";
					when "101100010011000" => rgb <= "101111";
					when "101100010011001" => rgb <= "101111";
					when "101100010011010" => rgb <= "101111";
					when "101100010011011" => rgb <= "101111";
					when "101100010011100" => rgb <= "101111";
					when "101100010011101" => rgb <= "101111";
					when "101100010011110" => rgb <= "101111";
					when "101100010011111" => rgb <= "101111";
					when "101100100000000" => rgb <= "101111";
					when "101100100000001" => rgb <= "101111";
					when "101100100000010" => rgb <= "101111";
					when "101100100000011" => rgb <= "101111";
					when "101100100000100" => rgb <= "101111";
					when "101100100000101" => rgb <= "101111";
					when "101100100000110" => rgb <= "101111";
					when "101100100000111" => rgb <= "101111";
					when "101100100001000" => rgb <= "101111";
					when "101100100001001" => rgb <= "101111";
					when "101100100001010" => rgb <= "101111";
					when "101100100001011" => rgb <= "101111";
					when "101100100001100" => rgb <= "101111";
					when "101100100001101" => rgb <= "101111";
					when "101100100001110" => rgb <= "101111";
					when "101100100001111" => rgb <= "101111";
					when "101100100010000" => rgb <= "101111";
					when "101100100010001" => rgb <= "101111";
					when "101100100010010" => rgb <= "101111";
					when "101100100010011" => rgb <= "101111";
					when "101100100010100" => rgb <= "101111";
					when "101100100010101" => rgb <= "101111";
					when "101100100010110" => rgb <= "101111";
					when "101100100010111" => rgb <= "101111";
					when "101100100011000" => rgb <= "101111";
					when "101100100011001" => rgb <= "101111";
					when "101100100011010" => rgb <= "101111";
					when "101100100011011" => rgb <= "101111";
					when "101100100011100" => rgb <= "101111";
					when "101100100011101" => rgb <= "101111";
					when "101100100011110" => rgb <= "101111";
					when "101100100011111" => rgb <= "101111";
					when "101100100100000" => rgb <= "000000";
					when "101100100100001" => rgb <= "000000";
					when "101100100100010" => rgb <= "100100";
					when "101100100100011" => rgb <= "100100";
					when "101100100100100" => rgb <= "100100";
					when "101100100100101" => rgb <= "100100";
					when "101100100100110" => rgb <= "100100";
					when "101100100100111" => rgb <= "100100";
					when "101100100101000" => rgb <= "100100";
					when "101100100101001" => rgb <= "100100";
					when "101100100101010" => rgb <= "100100";
					when "101100100101011" => rgb <= "100100";
					when "101100100101100" => rgb <= "100100";
					when "101100100101101" => rgb <= "100100";
					when "101100100101110" => rgb <= "100100";
					when "101100100101111" => rgb <= "100100";
					when "101100100110000" => rgb <= "100100";
					when "101100100110001" => rgb <= "100100";
					when "101100100110010" => rgb <= "010000";
					when "101100100110011" => rgb <= "010000";
					when "101100100110100" => rgb <= "000000";
					when "101100100110101" => rgb <= "000000";
					when "101100100110110" => rgb <= "101111";
					when "101100100110111" => rgb <= "101111";
					when "101100100111000" => rgb <= "101111";
					when "101100100111001" => rgb <= "101111";
					when "101100100111010" => rgb <= "101111";
					when "101100100111011" => rgb <= "101111";
					when "101100100111100" => rgb <= "101111";
					when "101100100111101" => rgb <= "101111";
					when "101100100111110" => rgb <= "101111";
					when "101100100111111" => rgb <= "101111";
					when "101100101000000" => rgb <= "101111";
					when "101100101000001" => rgb <= "101111";
					when "101100101000010" => rgb <= "101111";
					when "101100101000011" => rgb <= "101111";
					when "101100101000100" => rgb <= "101111";
					when "101100101000101" => rgb <= "101111";
					when "101100101000110" => rgb <= "101111";
					when "101100101000111" => rgb <= "101111";
					when "101100101001000" => rgb <= "101111";
					when "101100101001001" => rgb <= "101111";
					when "101100101001010" => rgb <= "101111";
					when "101100101001011" => rgb <= "101111";
					when "101100101001100" => rgb <= "101111";
					when "101100101001101" => rgb <= "101111";
					when "101100101001110" => rgb <= "101111";
					when "101100101001111" => rgb <= "101111";
					when "101100101010000" => rgb <= "101111";
					when "101100101010001" => rgb <= "101111";
					when "101100101010010" => rgb <= "101111";
					when "101100101010011" => rgb <= "101111";
					when "101100101010100" => rgb <= "101111";
					when "101100101010101" => rgb <= "101111";
					when "101100101010110" => rgb <= "101111";
					when "101100101010111" => rgb <= "101111";
					when "101100101011000" => rgb <= "101111";
					when "101100101011001" => rgb <= "101111";
					when "101100101011010" => rgb <= "101111";
					when "101100101011011" => rgb <= "101111";
					when "101100101011100" => rgb <= "101111";
					when "101100101011101" => rgb <= "101111";
					when "101100101011110" => rgb <= "101111";
					when "101100101011111" => rgb <= "101111";
					when "101100101100000" => rgb <= "101111";
					when "101100101100001" => rgb <= "101111";
					when "101100101100010" => rgb <= "101111";
					when "101100101100011" => rgb <= "101111";
					when "101100101100100" => rgb <= "101111";
					when "101100101100101" => rgb <= "101111";
					when "101100101100110" => rgb <= "101111";
					when "101100101100111" => rgb <= "101111";
					when "101100101101000" => rgb <= "101111";
					when "101100101101001" => rgb <= "101111";
					when "101100101101010" => rgb <= "101111";
					when "101100101101011" => rgb <= "101111";
					when "101100101101100" => rgb <= "101111";
					when "101100101101101" => rgb <= "101111";
					when "101100101101110" => rgb <= "101111";
					when "101100101101111" => rgb <= "101111";
					when "101100101110000" => rgb <= "101111";
					when "101100101110001" => rgb <= "101111";
					when "101100101110010" => rgb <= "101111";
					when "101100101110011" => rgb <= "101111";
					when "101100101110100" => rgb <= "101111";
					when "101100101110101" => rgb <= "101111";
					when "101100101110110" => rgb <= "101111";
					when "101100101110111" => rgb <= "101111";
					when "101100101111000" => rgb <= "101111";
					when "101100101111001" => rgb <= "101111";
					when "101100101111010" => rgb <= "101111";
					when "101100101111011" => rgb <= "101111";
					when "101100101111100" => rgb <= "101111";
					when "101100101111101" => rgb <= "101111";
					when "101100101111110" => rgb <= "101111";
					when "101100101111111" => rgb <= "101111";
					when "101100110000000" => rgb <= "101111";
					when "101100110000001" => rgb <= "101111";
					when "101100110000010" => rgb <= "101111";
					when "101100110000011" => rgb <= "101111";
					when "101100110000100" => rgb <= "101111";
					when "101100110000101" => rgb <= "101111";
					when "101100110000110" => rgb <= "101111";
					when "101100110000111" => rgb <= "101111";
					when "101100110001000" => rgb <= "101111";
					when "101100110001001" => rgb <= "101111";
					when "101100110001010" => rgb <= "101111";
					when "101100110001011" => rgb <= "101111";
					when "101100110001100" => rgb <= "101111";
					when "101100110001101" => rgb <= "101111";
					when "101100110001110" => rgb <= "101111";
					when "101100110001111" => rgb <= "101111";
					when "101100110010000" => rgb <= "101111";
					when "101100110010001" => rgb <= "101111";
					when "101100110010010" => rgb <= "101111";
					when "101100110010011" => rgb <= "101111";
					when "101100110010100" => rgb <= "101111";
					when "101100110010101" => rgb <= "101111";
					when "101100110010110" => rgb <= "101111";
					when "101100110010111" => rgb <= "101111";
					when "101100110011000" => rgb <= "101111";
					when "101100110011001" => rgb <= "101111";
					when "101100110011010" => rgb <= "101111";
					when "101100110011011" => rgb <= "101111";
					when "101100110011100" => rgb <= "101111";
					when "101100110011101" => rgb <= "101111";
					when "101100110011110" => rgb <= "101111";
					when "101100110011111" => rgb <= "101111";
					when "101101000000000" => rgb <= "101111";
					when "101101000000001" => rgb <= "101111";
					when "101101000000010" => rgb <= "101111";
					when "101101000000011" => rgb <= "101111";
					when "101101000000100" => rgb <= "101111";
					when "101101000000101" => rgb <= "101111";
					when "101101000000110" => rgb <= "101111";
					when "101101000000111" => rgb <= "101111";
					when "101101000001000" => rgb <= "101111";
					when "101101000001001" => rgb <= "101111";
					when "101101000001010" => rgb <= "101111";
					when "101101000001011" => rgb <= "101111";
					when "101101000001100" => rgb <= "101111";
					when "101101000001101" => rgb <= "101111";
					when "101101000001110" => rgb <= "101111";
					when "101101000001111" => rgb <= "101111";
					when "101101000010000" => rgb <= "101111";
					when "101101000010001" => rgb <= "101111";
					when "101101000010010" => rgb <= "101111";
					when "101101000010011" => rgb <= "101111";
					when "101101000010100" => rgb <= "101111";
					when "101101000010101" => rgb <= "101111";
					when "101101000010110" => rgb <= "101111";
					when "101101000010111" => rgb <= "101111";
					when "101101000011000" => rgb <= "101111";
					when "101101000011001" => rgb <= "101111";
					when "101101000011010" => rgb <= "101111";
					when "101101000011011" => rgb <= "101111";
					when "101101000011100" => rgb <= "101111";
					when "101101000011101" => rgb <= "101111";
					when "101101000011110" => rgb <= "101111";
					when "101101000011111" => rgb <= "101111";
					when "101101000100000" => rgb <= "000000";
					when "101101000100001" => rgb <= "000000";
					when "101101000100010" => rgb <= "100100";
					when "101101000100011" => rgb <= "100100";
					when "101101000100100" => rgb <= "100100";
					when "101101000100101" => rgb <= "100100";
					when "101101000100110" => rgb <= "100100";
					when "101101000100111" => rgb <= "100100";
					when "101101000101000" => rgb <= "100100";
					when "101101000101001" => rgb <= "100100";
					when "101101000101010" => rgb <= "100100";
					when "101101000101011" => rgb <= "100100";
					when "101101000101100" => rgb <= "100100";
					when "101101000101101" => rgb <= "100100";
					when "101101000101110" => rgb <= "100100";
					when "101101000101111" => rgb <= "100100";
					when "101101000110000" => rgb <= "100100";
					when "101101000110001" => rgb <= "100100";
					when "101101000110010" => rgb <= "010000";
					when "101101000110011" => rgb <= "010000";
					when "101101000110100" => rgb <= "000000";
					when "101101000110101" => rgb <= "000000";
					when "101101000110110" => rgb <= "101111";
					when "101101000110111" => rgb <= "101111";
					when "101101000111000" => rgb <= "101111";
					when "101101000111001" => rgb <= "101111";
					when "101101000111010" => rgb <= "101111";
					when "101101000111011" => rgb <= "101111";
					when "101101000111100" => rgb <= "101111";
					when "101101000111101" => rgb <= "101111";
					when "101101000111110" => rgb <= "101111";
					when "101101000111111" => rgb <= "101111";
					when "101101001000000" => rgb <= "101111";
					when "101101001000001" => rgb <= "101111";
					when "101101001000010" => rgb <= "101111";
					when "101101001000011" => rgb <= "101111";
					when "101101001000100" => rgb <= "101111";
					when "101101001000101" => rgb <= "101111";
					when "101101001000110" => rgb <= "101111";
					when "101101001000111" => rgb <= "101111";
					when "101101001001000" => rgb <= "101111";
					when "101101001001001" => rgb <= "101111";
					when "101101001001010" => rgb <= "101111";
					when "101101001001011" => rgb <= "101111";
					when "101101001001100" => rgb <= "101111";
					when "101101001001101" => rgb <= "101111";
					when "101101001001110" => rgb <= "101111";
					when "101101001001111" => rgb <= "101111";
					when "101101001010000" => rgb <= "101111";
					when "101101001010001" => rgb <= "101111";
					when "101101001010010" => rgb <= "101111";
					when "101101001010011" => rgb <= "101111";
					when "101101001010100" => rgb <= "101111";
					when "101101001010101" => rgb <= "101111";
					when "101101001010110" => rgb <= "101111";
					when "101101001010111" => rgb <= "101111";
					when "101101001011000" => rgb <= "101111";
					when "101101001011001" => rgb <= "101111";
					when "101101001011010" => rgb <= "101111";
					when "101101001011011" => rgb <= "101111";
					when "101101001011100" => rgb <= "101111";
					when "101101001011101" => rgb <= "101111";
					when "101101001011110" => rgb <= "101111";
					when "101101001011111" => rgb <= "101111";
					when "101101001100000" => rgb <= "101111";
					when "101101001100001" => rgb <= "101111";
					when "101101001100010" => rgb <= "101111";
					when "101101001100011" => rgb <= "101111";
					when "101101001100100" => rgb <= "101111";
					when "101101001100101" => rgb <= "101111";
					when "101101001100110" => rgb <= "101111";
					when "101101001100111" => rgb <= "101111";
					when "101101001101000" => rgb <= "101111";
					when "101101001101001" => rgb <= "101111";
					when "101101001101010" => rgb <= "101111";
					when "101101001101011" => rgb <= "101111";
					when "101101001101100" => rgb <= "101111";
					when "101101001101101" => rgb <= "101111";
					when "101101001101110" => rgb <= "101111";
					when "101101001101111" => rgb <= "101111";
					when "101101001110000" => rgb <= "101111";
					when "101101001110001" => rgb <= "101111";
					when "101101001110010" => rgb <= "101111";
					when "101101001110011" => rgb <= "101111";
					when "101101001110100" => rgb <= "101111";
					when "101101001110101" => rgb <= "101111";
					when "101101001110110" => rgb <= "101111";
					when "101101001110111" => rgb <= "101111";
					when "101101001111000" => rgb <= "101111";
					when "101101001111001" => rgb <= "101111";
					when "101101001111010" => rgb <= "101111";
					when "101101001111011" => rgb <= "101111";
					when "101101001111100" => rgb <= "101111";
					when "101101001111101" => rgb <= "101111";
					when "101101001111110" => rgb <= "101111";
					when "101101001111111" => rgb <= "101111";
					when "101101010000000" => rgb <= "101111";
					when "101101010000001" => rgb <= "101111";
					when "101101010000010" => rgb <= "101111";
					when "101101010000011" => rgb <= "101111";
					when "101101010000100" => rgb <= "101111";
					when "101101010000101" => rgb <= "101111";
					when "101101010000110" => rgb <= "101111";
					when "101101010000111" => rgb <= "101111";
					when "101101010001000" => rgb <= "101111";
					when "101101010001001" => rgb <= "101111";
					when "101101010001010" => rgb <= "101111";
					when "101101010001011" => rgb <= "101111";
					when "101101010001100" => rgb <= "101111";
					when "101101010001101" => rgb <= "101111";
					when "101101010001110" => rgb <= "101111";
					when "101101010001111" => rgb <= "101111";
					when "101101010010000" => rgb <= "101111";
					when "101101010010001" => rgb <= "101111";
					when "101101010010010" => rgb <= "101111";
					when "101101010010011" => rgb <= "101111";
					when "101101010010100" => rgb <= "101111";
					when "101101010010101" => rgb <= "101111";
					when "101101010010110" => rgb <= "101111";
					when "101101010010111" => rgb <= "101111";
					when "101101010011000" => rgb <= "101111";
					when "101101010011001" => rgb <= "101111";
					when "101101010011010" => rgb <= "101111";
					when "101101010011011" => rgb <= "101111";
					when "101101010011100" => rgb <= "101111";
					when "101101010011101" => rgb <= "101111";
					when "101101010011110" => rgb <= "101111";
					when "101101010011111" => rgb <= "101111";
					when "101101100000000" => rgb <= "101111";
					when "101101100000001" => rgb <= "101111";
					when "101101100000010" => rgb <= "101111";
					when "101101100000011" => rgb <= "101111";
					when "101101100000100" => rgb <= "101111";
					when "101101100000101" => rgb <= "101111";
					when "101101100000110" => rgb <= "101111";
					when "101101100000111" => rgb <= "101111";
					when "101101100001000" => rgb <= "101111";
					when "101101100001001" => rgb <= "101111";
					when "101101100001010" => rgb <= "101111";
					when "101101100001011" => rgb <= "101111";
					when "101101100001100" => rgb <= "101111";
					when "101101100001101" => rgb <= "101111";
					when "101101100001110" => rgb <= "101111";
					when "101101100001111" => rgb <= "101111";
					when "101101100010000" => rgb <= "101111";
					when "101101100010001" => rgb <= "101111";
					when "101101100010010" => rgb <= "101111";
					when "101101100010011" => rgb <= "101111";
					when "101101100010100" => rgb <= "101111";
					when "101101100010101" => rgb <= "101111";
					when "101101100010110" => rgb <= "101111";
					when "101101100010111" => rgb <= "101111";
					when "101101100011000" => rgb <= "101111";
					when "101101100011001" => rgb <= "101111";
					when "101101100011010" => rgb <= "101111";
					when "101101100011011" => rgb <= "101111";
					when "101101100011100" => rgb <= "101111";
					when "101101100011101" => rgb <= "101111";
					when "101101100011110" => rgb <= "101111";
					when "101101100011111" => rgb <= "101111";
					when "101101100100000" => rgb <= "000000";
					when "101101100100001" => rgb <= "000000";
					when "101101100100010" => rgb <= "100100";
					when "101101100100011" => rgb <= "100100";
					when "101101100100100" => rgb <= "100100";
					when "101101100100101" => rgb <= "100100";
					when "101101100100110" => rgb <= "100100";
					when "101101100100111" => rgb <= "100100";
					when "101101100101000" => rgb <= "100100";
					when "101101100101001" => rgb <= "100100";
					when "101101100101010" => rgb <= "100100";
					when "101101100101011" => rgb <= "100100";
					when "101101100101100" => rgb <= "100100";
					when "101101100101101" => rgb <= "100100";
					when "101101100101110" => rgb <= "100100";
					when "101101100101111" => rgb <= "100100";
					when "101101100110000" => rgb <= "100100";
					when "101101100110001" => rgb <= "100100";
					when "101101100110010" => rgb <= "010000";
					when "101101100110011" => rgb <= "010000";
					when "101101100110100" => rgb <= "000000";
					when "101101100110101" => rgb <= "000000";
					when "101101100110110" => rgb <= "101111";
					when "101101100110111" => rgb <= "101111";
					when "101101100111000" => rgb <= "101111";
					when "101101100111001" => rgb <= "101111";
					when "101101100111010" => rgb <= "101111";
					when "101101100111011" => rgb <= "101111";
					when "101101100111100" => rgb <= "101111";
					when "101101100111101" => rgb <= "101111";
					when "101101100111110" => rgb <= "101111";
					when "101101100111111" => rgb <= "101111";
					when "101101101000000" => rgb <= "101111";
					when "101101101000001" => rgb <= "101111";
					when "101101101000010" => rgb <= "101111";
					when "101101101000011" => rgb <= "101111";
					when "101101101000100" => rgb <= "101111";
					when "101101101000101" => rgb <= "101111";
					when "101101101000110" => rgb <= "101111";
					when "101101101000111" => rgb <= "101111";
					when "101101101001000" => rgb <= "101111";
					when "101101101001001" => rgb <= "101111";
					when "101101101001010" => rgb <= "101111";
					when "101101101001011" => rgb <= "101111";
					when "101101101001100" => rgb <= "101111";
					when "101101101001101" => rgb <= "101111";
					when "101101101001110" => rgb <= "101111";
					when "101101101001111" => rgb <= "101111";
					when "101101101010000" => rgb <= "101111";
					when "101101101010001" => rgb <= "101111";
					when "101101101010010" => rgb <= "101111";
					when "101101101010011" => rgb <= "101111";
					when "101101101010100" => rgb <= "101111";
					when "101101101010101" => rgb <= "101111";
					when "101101101010110" => rgb <= "101111";
					when "101101101010111" => rgb <= "101111";
					when "101101101011000" => rgb <= "101111";
					when "101101101011001" => rgb <= "101111";
					when "101101101011010" => rgb <= "101111";
					when "101101101011011" => rgb <= "101111";
					when "101101101011100" => rgb <= "101111";
					when "101101101011101" => rgb <= "101111";
					when "101101101011110" => rgb <= "101111";
					when "101101101011111" => rgb <= "101111";
					when "101101101100000" => rgb <= "101111";
					when "101101101100001" => rgb <= "101111";
					when "101101101100010" => rgb <= "101111";
					when "101101101100011" => rgb <= "101111";
					when "101101101100100" => rgb <= "101111";
					when "101101101100101" => rgb <= "101111";
					when "101101101100110" => rgb <= "101111";
					when "101101101100111" => rgb <= "101111";
					when "101101101101000" => rgb <= "101111";
					when "101101101101001" => rgb <= "101111";
					when "101101101101010" => rgb <= "101111";
					when "101101101101011" => rgb <= "101111";
					when "101101101101100" => rgb <= "101111";
					when "101101101101101" => rgb <= "101111";
					when "101101101101110" => rgb <= "101111";
					when "101101101101111" => rgb <= "101111";
					when "101101101110000" => rgb <= "101111";
					when "101101101110001" => rgb <= "101111";
					when "101101101110010" => rgb <= "101111";
					when "101101101110011" => rgb <= "101111";
					when "101101101110100" => rgb <= "101111";
					when "101101101110101" => rgb <= "101111";
					when "101101101110110" => rgb <= "101111";
					when "101101101110111" => rgb <= "101111";
					when "101101101111000" => rgb <= "101111";
					when "101101101111001" => rgb <= "101111";
					when "101101101111010" => rgb <= "101111";
					when "101101101111011" => rgb <= "101111";
					when "101101101111100" => rgb <= "101111";
					when "101101101111101" => rgb <= "101111";
					when "101101101111110" => rgb <= "101111";
					when "101101101111111" => rgb <= "101111";
					when "101101110000000" => rgb <= "101111";
					when "101101110000001" => rgb <= "101111";
					when "101101110000010" => rgb <= "101111";
					when "101101110000011" => rgb <= "101111";
					when "101101110000100" => rgb <= "101111";
					when "101101110000101" => rgb <= "101111";
					when "101101110000110" => rgb <= "101111";
					when "101101110000111" => rgb <= "101111";
					when "101101110001000" => rgb <= "101111";
					when "101101110001001" => rgb <= "101111";
					when "101101110001010" => rgb <= "101111";
					when "101101110001011" => rgb <= "101111";
					when "101101110001100" => rgb <= "101111";
					when "101101110001101" => rgb <= "101111";
					when "101101110001110" => rgb <= "101111";
					when "101101110001111" => rgb <= "101111";
					when "101101110010000" => rgb <= "101111";
					when "101101110010001" => rgb <= "101111";
					when "101101110010010" => rgb <= "101111";
					when "101101110010011" => rgb <= "101111";
					when "101101110010100" => rgb <= "101111";
					when "101101110010101" => rgb <= "101111";
					when "101101110010110" => rgb <= "101111";
					when "101101110010111" => rgb <= "101111";
					when "101101110011000" => rgb <= "101111";
					when "101101110011001" => rgb <= "101111";
					when "101101110011010" => rgb <= "101111";
					when "101101110011011" => rgb <= "101111";
					when "101101110011100" => rgb <= "101111";
					when "101101110011101" => rgb <= "101111";
					when "101101110011110" => rgb <= "101111";
					when "101101110011111" => rgb <= "101111";
					when "101110000000000" => rgb <= "101111";
					when "101110000000001" => rgb <= "101111";
					when "101110000000010" => rgb <= "101111";
					when "101110000000011" => rgb <= "101111";
					when "101110000000100" => rgb <= "101111";
					when "101110000000101" => rgb <= "101111";
					when "101110000000110" => rgb <= "101111";
					when "101110000000111" => rgb <= "101111";
					when "101110000001000" => rgb <= "101111";
					when "101110000001001" => rgb <= "101111";
					when "101110000001010" => rgb <= "101111";
					when "101110000001011" => rgb <= "101111";
					when "101110000001100" => rgb <= "101111";
					when "101110000001101" => rgb <= "101111";
					when "101110000001110" => rgb <= "101111";
					when "101110000001111" => rgb <= "101111";
					when "101110000010000" => rgb <= "101111";
					when "101110000010001" => rgb <= "101111";
					when "101110000010010" => rgb <= "101111";
					when "101110000010011" => rgb <= "101111";
					when "101110000010100" => rgb <= "101111";
					when "101110000010101" => rgb <= "101111";
					when "101110000010110" => rgb <= "101111";
					when "101110000010111" => rgb <= "101111";
					when "101110000011000" => rgb <= "101111";
					when "101110000011001" => rgb <= "101111";
					when "101110000011010" => rgb <= "101111";
					when "101110000011011" => rgb <= "101111";
					when "101110000011100" => rgb <= "101111";
					when "101110000011101" => rgb <= "101111";
					when "101110000011110" => rgb <= "101111";
					when "101110000011111" => rgb <= "101111";
					when "101110000100000" => rgb <= "000000";
					when "101110000100001" => rgb <= "000000";
					when "101110000100010" => rgb <= "100100";
					when "101110000100011" => rgb <= "100100";
					when "101110000100100" => rgb <= "100100";
					when "101110000100101" => rgb <= "100100";
					when "101110000100110" => rgb <= "100100";
					when "101110000100111" => rgb <= "100100";
					when "101110000101000" => rgb <= "100100";
					when "101110000101001" => rgb <= "100100";
					when "101110000101010" => rgb <= "100100";
					when "101110000101011" => rgb <= "100100";
					when "101110000101100" => rgb <= "100100";
					when "101110000101101" => rgb <= "100100";
					when "101110000101110" => rgb <= "100100";
					when "101110000101111" => rgb <= "100100";
					when "101110000110000" => rgb <= "100100";
					when "101110000110001" => rgb <= "100100";
					when "101110000110010" => rgb <= "010000";
					when "101110000110011" => rgb <= "010000";
					when "101110000110100" => rgb <= "000000";
					when "101110000110101" => rgb <= "000000";
					when "101110000110110" => rgb <= "101111";
					when "101110000110111" => rgb <= "101111";
					when "101110000111000" => rgb <= "101111";
					when "101110000111001" => rgb <= "101111";
					when "101110000111010" => rgb <= "101111";
					when "101110000111011" => rgb <= "101111";
					when "101110000111100" => rgb <= "101111";
					when "101110000111101" => rgb <= "101111";
					when "101110000111110" => rgb <= "101111";
					when "101110000111111" => rgb <= "101111";
					when "101110001000000" => rgb <= "101111";
					when "101110001000001" => rgb <= "101111";
					when "101110001000010" => rgb <= "101111";
					when "101110001000011" => rgb <= "101111";
					when "101110001000100" => rgb <= "101111";
					when "101110001000101" => rgb <= "101111";
					when "101110001000110" => rgb <= "101111";
					when "101110001000111" => rgb <= "101111";
					when "101110001001000" => rgb <= "101111";
					when "101110001001001" => rgb <= "101111";
					when "101110001001010" => rgb <= "101111";
					when "101110001001011" => rgb <= "101111";
					when "101110001001100" => rgb <= "101111";
					when "101110001001101" => rgb <= "101111";
					when "101110001001110" => rgb <= "101111";
					when "101110001001111" => rgb <= "101111";
					when "101110001010000" => rgb <= "101111";
					when "101110001010001" => rgb <= "101111";
					when "101110001010010" => rgb <= "101111";
					when "101110001010011" => rgb <= "101111";
					when "101110001010100" => rgb <= "101111";
					when "101110001010101" => rgb <= "101111";
					when "101110001010110" => rgb <= "101111";
					when "101110001010111" => rgb <= "101111";
					when "101110001011000" => rgb <= "101111";
					when "101110001011001" => rgb <= "101111";
					when "101110001011010" => rgb <= "101111";
					when "101110001011011" => rgb <= "101111";
					when "101110001011100" => rgb <= "101111";
					when "101110001011101" => rgb <= "101111";
					when "101110001011110" => rgb <= "101111";
					when "101110001011111" => rgb <= "101111";
					when "101110001100000" => rgb <= "101111";
					when "101110001100001" => rgb <= "101111";
					when "101110001100010" => rgb <= "101111";
					when "101110001100011" => rgb <= "101111";
					when "101110001100100" => rgb <= "101111";
					when "101110001100101" => rgb <= "101111";
					when "101110001100110" => rgb <= "101111";
					when "101110001100111" => rgb <= "101111";
					when "101110001101000" => rgb <= "101111";
					when "101110001101001" => rgb <= "101111";
					when "101110001101010" => rgb <= "101111";
					when "101110001101011" => rgb <= "101111";
					when "101110001101100" => rgb <= "101111";
					when "101110001101101" => rgb <= "101111";
					when "101110001101110" => rgb <= "101111";
					when "101110001101111" => rgb <= "101111";
					when "101110001110000" => rgb <= "101111";
					when "101110001110001" => rgb <= "101111";
					when "101110001110010" => rgb <= "101111";
					when "101110001110011" => rgb <= "101111";
					when "101110001110100" => rgb <= "101111";
					when "101110001110101" => rgb <= "101111";
					when "101110001110110" => rgb <= "101111";
					when "101110001110111" => rgb <= "101111";
					when "101110001111000" => rgb <= "101111";
					when "101110001111001" => rgb <= "101111";
					when "101110001111010" => rgb <= "101111";
					when "101110001111011" => rgb <= "101111";
					when "101110001111100" => rgb <= "101111";
					when "101110001111101" => rgb <= "101111";
					when "101110001111110" => rgb <= "101111";
					when "101110001111111" => rgb <= "101111";
					when "101110010000000" => rgb <= "101111";
					when "101110010000001" => rgb <= "101111";
					when "101110010000010" => rgb <= "101111";
					when "101110010000011" => rgb <= "101111";
					when "101110010000100" => rgb <= "101111";
					when "101110010000101" => rgb <= "101111";
					when "101110010000110" => rgb <= "101111";
					when "101110010000111" => rgb <= "101111";
					when "101110010001000" => rgb <= "101111";
					when "101110010001001" => rgb <= "101111";
					when "101110010001010" => rgb <= "101111";
					when "101110010001011" => rgb <= "101111";
					when "101110010001100" => rgb <= "101111";
					when "101110010001101" => rgb <= "101111";
					when "101110010001110" => rgb <= "101111";
					when "101110010001111" => rgb <= "101111";
					when "101110010010000" => rgb <= "101111";
					when "101110010010001" => rgb <= "101111";
					when "101110010010010" => rgb <= "101111";
					when "101110010010011" => rgb <= "101111";
					when "101110010010100" => rgb <= "101111";
					when "101110010010101" => rgb <= "101111";
					when "101110010010110" => rgb <= "101111";
					when "101110010010111" => rgb <= "101111";
					when "101110010011000" => rgb <= "101111";
					when "101110010011001" => rgb <= "101111";
					when "101110010011010" => rgb <= "101111";
					when "101110010011011" => rgb <= "101111";
					when "101110010011100" => rgb <= "101111";
					when "101110010011101" => rgb <= "101111";
					when "101110010011110" => rgb <= "101111";
					when "101110010011111" => rgb <= "101111";
					when "101110100000000" => rgb <= "101111";
					when "101110100000001" => rgb <= "101111";
					when "101110100000010" => rgb <= "101111";
					when "101110100000011" => rgb <= "101111";
					when "101110100000100" => rgb <= "101111";
					when "101110100000101" => rgb <= "101111";
					when "101110100000110" => rgb <= "101111";
					when "101110100000111" => rgb <= "101111";
					when "101110100001000" => rgb <= "101111";
					when "101110100001001" => rgb <= "101111";
					when "101110100001010" => rgb <= "101111";
					when "101110100001011" => rgb <= "101111";
					when "101110100001100" => rgb <= "101111";
					when "101110100001101" => rgb <= "101111";
					when "101110100001110" => rgb <= "101111";
					when "101110100001111" => rgb <= "101111";
					when "101110100010000" => rgb <= "101111";
					when "101110100010001" => rgb <= "101111";
					when "101110100010010" => rgb <= "101111";
					when "101110100010011" => rgb <= "101111";
					when "101110100010100" => rgb <= "101111";
					when "101110100010101" => rgb <= "101111";
					when "101110100010110" => rgb <= "101111";
					when "101110100010111" => rgb <= "101111";
					when "101110100011000" => rgb <= "101111";
					when "101110100011001" => rgb <= "101111";
					when "101110100011010" => rgb <= "101111";
					when "101110100011011" => rgb <= "101111";
					when "101110100011100" => rgb <= "101111";
					when "101110100011101" => rgb <= "101111";
					when "101110100011110" => rgb <= "101111";
					when "101110100011111" => rgb <= "101111";
					when "101110100100000" => rgb <= "000000";
					when "101110100100001" => rgb <= "000000";
					when "101110100100010" => rgb <= "100100";
					when "101110100100011" => rgb <= "100100";
					when "101110100100100" => rgb <= "100100";
					when "101110100100101" => rgb <= "100100";
					when "101110100100110" => rgb <= "100100";
					when "101110100100111" => rgb <= "100100";
					when "101110100101000" => rgb <= "100100";
					when "101110100101001" => rgb <= "100100";
					when "101110100101010" => rgb <= "100100";
					when "101110100101011" => rgb <= "100100";
					when "101110100101100" => rgb <= "100100";
					when "101110100101101" => rgb <= "100100";
					when "101110100101110" => rgb <= "100100";
					when "101110100101111" => rgb <= "100100";
					when "101110100110000" => rgb <= "100100";
					when "101110100110001" => rgb <= "100100";
					when "101110100110010" => rgb <= "010000";
					when "101110100110011" => rgb <= "010000";
					when "101110100110100" => rgb <= "000000";
					when "101110100110101" => rgb <= "000000";
					when "101110100110110" => rgb <= "101111";
					when "101110100110111" => rgb <= "101111";
					when "101110100111000" => rgb <= "101111";
					when "101110100111001" => rgb <= "101111";
					when "101110100111010" => rgb <= "101111";
					when "101110100111011" => rgb <= "101111";
					when "101110100111100" => rgb <= "101111";
					when "101110100111101" => rgb <= "101111";
					when "101110100111110" => rgb <= "101111";
					when "101110100111111" => rgb <= "101111";
					when "101110101000000" => rgb <= "101111";
					when "101110101000001" => rgb <= "101111";
					when "101110101000010" => rgb <= "101111";
					when "101110101000011" => rgb <= "101111";
					when "101110101000100" => rgb <= "101111";
					when "101110101000101" => rgb <= "101111";
					when "101110101000110" => rgb <= "101111";
					when "101110101000111" => rgb <= "101111";
					when "101110101001000" => rgb <= "101111";
					when "101110101001001" => rgb <= "101111";
					when "101110101001010" => rgb <= "101111";
					when "101110101001011" => rgb <= "101111";
					when "101110101001100" => rgb <= "101111";
					when "101110101001101" => rgb <= "101111";
					when "101110101001110" => rgb <= "101111";
					when "101110101001111" => rgb <= "101111";
					when "101110101010000" => rgb <= "101111";
					when "101110101010001" => rgb <= "101111";
					when "101110101010010" => rgb <= "101111";
					when "101110101010011" => rgb <= "101111";
					when "101110101010100" => rgb <= "101111";
					when "101110101010101" => rgb <= "101111";
					when "101110101010110" => rgb <= "101111";
					when "101110101010111" => rgb <= "101111";
					when "101110101011000" => rgb <= "101111";
					when "101110101011001" => rgb <= "101111";
					when "101110101011010" => rgb <= "101111";
					when "101110101011011" => rgb <= "101111";
					when "101110101011100" => rgb <= "101111";
					when "101110101011101" => rgb <= "101111";
					when "101110101011110" => rgb <= "101111";
					when "101110101011111" => rgb <= "101111";
					when "101110101100000" => rgb <= "101111";
					when "101110101100001" => rgb <= "101111";
					when "101110101100010" => rgb <= "101111";
					when "101110101100011" => rgb <= "101111";
					when "101110101100100" => rgb <= "101111";
					when "101110101100101" => rgb <= "101111";
					when "101110101100110" => rgb <= "101111";
					when "101110101100111" => rgb <= "101111";
					when "101110101101000" => rgb <= "101111";
					when "101110101101001" => rgb <= "101111";
					when "101110101101010" => rgb <= "101111";
					when "101110101101011" => rgb <= "101111";
					when "101110101101100" => rgb <= "101111";
					when "101110101101101" => rgb <= "101111";
					when "101110101101110" => rgb <= "101111";
					when "101110101101111" => rgb <= "101111";
					when "101110101110000" => rgb <= "101111";
					when "101110101110001" => rgb <= "101111";
					when "101110101110010" => rgb <= "101111";
					when "101110101110011" => rgb <= "101111";
					when "101110101110100" => rgb <= "101111";
					when "101110101110101" => rgb <= "101111";
					when "101110101110110" => rgb <= "101111";
					when "101110101110111" => rgb <= "101111";
					when "101110101111000" => rgb <= "101111";
					when "101110101111001" => rgb <= "101111";
					when "101110101111010" => rgb <= "101111";
					when "101110101111011" => rgb <= "101111";
					when "101110101111100" => rgb <= "101111";
					when "101110101111101" => rgb <= "101111";
					when "101110101111110" => rgb <= "101111";
					when "101110101111111" => rgb <= "101111";
					when "101110110000000" => rgb <= "101111";
					when "101110110000001" => rgb <= "101111";
					when "101110110000010" => rgb <= "101111";
					when "101110110000011" => rgb <= "101111";
					when "101110110000100" => rgb <= "101111";
					when "101110110000101" => rgb <= "101111";
					when "101110110000110" => rgb <= "101111";
					when "101110110000111" => rgb <= "101111";
					when "101110110001000" => rgb <= "101111";
					when "101110110001001" => rgb <= "101111";
					when "101110110001010" => rgb <= "101111";
					when "101110110001011" => rgb <= "101111";
					when "101110110001100" => rgb <= "101111";
					when "101110110001101" => rgb <= "101111";
					when "101110110001110" => rgb <= "101111";
					when "101110110001111" => rgb <= "101111";
					when "101110110010000" => rgb <= "101111";
					when "101110110010001" => rgb <= "101111";
					when "101110110010010" => rgb <= "101111";
					when "101110110010011" => rgb <= "101111";
					when "101110110010100" => rgb <= "101111";
					when "101110110010101" => rgb <= "101111";
					when "101110110010110" => rgb <= "101111";
					when "101110110010111" => rgb <= "101111";
					when "101110110011000" => rgb <= "101111";
					when "101110110011001" => rgb <= "101111";
					when "101110110011010" => rgb <= "101111";
					when "101110110011011" => rgb <= "101111";
					when "101110110011100" => rgb <= "101111";
					when "101110110011101" => rgb <= "101111";
					when "101110110011110" => rgb <= "101111";
					when "101110110011111" => rgb <= "101111";
					when "101111000000000" => rgb <= "101111";
					when "101111000000001" => rgb <= "101111";
					when "101111000000010" => rgb <= "101111";
					when "101111000000011" => rgb <= "101111";
					when "101111000000100" => rgb <= "101111";
					when "101111000000101" => rgb <= "101111";
					when "101111000000110" => rgb <= "101111";
					when "101111000000111" => rgb <= "101111";
					when "101111000001000" => rgb <= "101111";
					when "101111000001001" => rgb <= "101111";
					when "101111000001010" => rgb <= "101111";
					when "101111000001011" => rgb <= "101111";
					when "101111000001100" => rgb <= "101111";
					when "101111000001101" => rgb <= "101111";
					when "101111000001110" => rgb <= "101111";
					when "101111000001111" => rgb <= "101111";
					when "101111000010000" => rgb <= "101111";
					when "101111000010001" => rgb <= "101111";
					when "101111000010010" => rgb <= "101111";
					when "101111000010011" => rgb <= "101111";
					when "101111000010100" => rgb <= "101111";
					when "101111000010101" => rgb <= "101111";
					when "101111000010110" => rgb <= "101111";
					when "101111000010111" => rgb <= "101111";
					when "101111000011000" => rgb <= "101111";
					when "101111000011001" => rgb <= "101111";
					when "101111000011010" => rgb <= "101111";
					when "101111000011011" => rgb <= "101111";
					when "101111000011100" => rgb <= "101111";
					when "101111000011101" => rgb <= "101111";
					when "101111000011110" => rgb <= "101111";
					when "101111000011111" => rgb <= "101111";
					when "101111000100000" => rgb <= "000000";
					when "101111000100001" => rgb <= "000000";
					when "101111000100010" => rgb <= "100100";
					when "101111000100011" => rgb <= "100100";
					when "101111000100100" => rgb <= "100100";
					when "101111000100101" => rgb <= "100100";
					when "101111000100110" => rgb <= "100100";
					when "101111000100111" => rgb <= "100100";
					when "101111000101000" => rgb <= "100100";
					when "101111000101001" => rgb <= "100100";
					when "101111000101010" => rgb <= "100100";
					when "101111000101011" => rgb <= "100100";
					when "101111000101100" => rgb <= "100100";
					when "101111000101101" => rgb <= "100100";
					when "101111000101110" => rgb <= "100100";
					when "101111000101111" => rgb <= "100100";
					when "101111000110000" => rgb <= "100100";
					when "101111000110001" => rgb <= "100100";
					when "101111000110010" => rgb <= "010000";
					when "101111000110011" => rgb <= "010000";
					when "101111000110100" => rgb <= "000000";
					when "101111000110101" => rgb <= "000000";
					when "101111000110110" => rgb <= "101111";
					when "101111000110111" => rgb <= "101111";
					when "101111000111000" => rgb <= "101111";
					when "101111000111001" => rgb <= "101111";
					when "101111000111010" => rgb <= "101111";
					when "101111000111011" => rgb <= "101111";
					when "101111000111100" => rgb <= "101111";
					when "101111000111101" => rgb <= "101111";
					when "101111000111110" => rgb <= "101111";
					when "101111000111111" => rgb <= "101111";
					when "101111001000000" => rgb <= "101111";
					when "101111001000001" => rgb <= "101111";
					when "101111001000010" => rgb <= "101111";
					when "101111001000011" => rgb <= "101111";
					when "101111001000100" => rgb <= "101111";
					when "101111001000101" => rgb <= "101111";
					when "101111001000110" => rgb <= "101111";
					when "101111001000111" => rgb <= "101111";
					when "101111001001000" => rgb <= "101111";
					when "101111001001001" => rgb <= "101111";
					when "101111001001010" => rgb <= "101111";
					when "101111001001011" => rgb <= "101111";
					when "101111001001100" => rgb <= "101111";
					when "101111001001101" => rgb <= "101111";
					when "101111001001110" => rgb <= "101111";
					when "101111001001111" => rgb <= "101111";
					when "101111001010000" => rgb <= "101111";
					when "101111001010001" => rgb <= "101111";
					when "101111001010010" => rgb <= "101111";
					when "101111001010011" => rgb <= "101111";
					when "101111001010100" => rgb <= "101111";
					when "101111001010101" => rgb <= "101111";
					when "101111001010110" => rgb <= "101111";
					when "101111001010111" => rgb <= "101111";
					when "101111001011000" => rgb <= "101111";
					when "101111001011001" => rgb <= "101111";
					when "101111001011010" => rgb <= "101111";
					when "101111001011011" => rgb <= "101111";
					when "101111001011100" => rgb <= "101111";
					when "101111001011101" => rgb <= "101111";
					when "101111001011110" => rgb <= "101111";
					when "101111001011111" => rgb <= "101111";
					when "101111001100000" => rgb <= "101111";
					when "101111001100001" => rgb <= "101111";
					when "101111001100010" => rgb <= "101111";
					when "101111001100011" => rgb <= "101111";
					when "101111001100100" => rgb <= "101111";
					when "101111001100101" => rgb <= "101111";
					when "101111001100110" => rgb <= "101111";
					when "101111001100111" => rgb <= "101111";
					when "101111001101000" => rgb <= "101111";
					when "101111001101001" => rgb <= "101111";
					when "101111001101010" => rgb <= "101111";
					when "101111001101011" => rgb <= "101111";
					when "101111001101100" => rgb <= "101111";
					when "101111001101101" => rgb <= "101111";
					when "101111001101110" => rgb <= "101111";
					when "101111001101111" => rgb <= "101111";
					when "101111001110000" => rgb <= "101111";
					when "101111001110001" => rgb <= "101111";
					when "101111001110010" => rgb <= "101111";
					when "101111001110011" => rgb <= "101111";
					when "101111001110100" => rgb <= "101111";
					when "101111001110101" => rgb <= "101111";
					when "101111001110110" => rgb <= "101111";
					when "101111001110111" => rgb <= "101111";
					when "101111001111000" => rgb <= "101111";
					when "101111001111001" => rgb <= "101111";
					when "101111001111010" => rgb <= "101111";
					when "101111001111011" => rgb <= "101111";
					when "101111001111100" => rgb <= "101111";
					when "101111001111101" => rgb <= "101111";
					when "101111001111110" => rgb <= "101111";
					when "101111001111111" => rgb <= "101111";
					when "101111010000000" => rgb <= "101111";
					when "101111010000001" => rgb <= "101111";
					when "101111010000010" => rgb <= "101111";
					when "101111010000011" => rgb <= "101111";
					when "101111010000100" => rgb <= "101111";
					when "101111010000101" => rgb <= "101111";
					when "101111010000110" => rgb <= "101111";
					when "101111010000111" => rgb <= "101111";
					when "101111010001000" => rgb <= "101111";
					when "101111010001001" => rgb <= "101111";
					when "101111010001010" => rgb <= "101111";
					when "101111010001011" => rgb <= "101111";
					when "101111010001100" => rgb <= "101111";
					when "101111010001101" => rgb <= "101111";
					when "101111010001110" => rgb <= "101111";
					when "101111010001111" => rgb <= "101111";
					when "101111010010000" => rgb <= "101111";
					when "101111010010001" => rgb <= "101111";
					when "101111010010010" => rgb <= "101111";
					when "101111010010011" => rgb <= "101111";
					when "101111010010100" => rgb <= "101111";
					when "101111010010101" => rgb <= "101111";
					when "101111010010110" => rgb <= "101111";
					when "101111010010111" => rgb <= "101111";
					when "101111010011000" => rgb <= "101111";
					when "101111010011001" => rgb <= "101111";
					when "101111010011010" => rgb <= "101111";
					when "101111010011011" => rgb <= "101111";
					when "101111010011100" => rgb <= "101111";
					when "101111010011101" => rgb <= "101111";
					when "101111010011110" => rgb <= "101111";
					when "101111010011111" => rgb <= "101111";
					when "101111100000000" => rgb <= "101111";
					when "101111100000001" => rgb <= "101111";
					when "101111100000010" => rgb <= "101111";
					when "101111100000011" => rgb <= "101111";
					when "101111100000100" => rgb <= "101111";
					when "101111100000101" => rgb <= "101111";
					when "101111100000110" => rgb <= "101111";
					when "101111100000111" => rgb <= "101111";
					when "101111100001000" => rgb <= "101111";
					when "101111100001001" => rgb <= "101111";
					when "101111100001010" => rgb <= "101111";
					when "101111100001011" => rgb <= "101111";
					when "101111100001100" => rgb <= "101111";
					when "101111100001101" => rgb <= "101111";
					when "101111100001110" => rgb <= "101111";
					when "101111100001111" => rgb <= "101111";
					when "101111100010000" => rgb <= "101111";
					when "101111100010001" => rgb <= "101111";
					when "101111100010010" => rgb <= "101111";
					when "101111100010011" => rgb <= "101111";
					when "101111100010100" => rgb <= "101111";
					when "101111100010101" => rgb <= "101111";
					when "101111100010110" => rgb <= "101111";
					when "101111100010111" => rgb <= "101111";
					when "101111100011000" => rgb <= "101111";
					when "101111100011001" => rgb <= "101111";
					when "101111100011010" => rgb <= "101111";
					when "101111100011011" => rgb <= "101111";
					when "101111100011100" => rgb <= "101111";
					when "101111100011101" => rgb <= "101111";
					when "101111100011110" => rgb <= "101111";
					when "101111100011111" => rgb <= "101111";
					when "101111100100000" => rgb <= "000000";
					when "101111100100001" => rgb <= "000000";
					when "101111100100010" => rgb <= "100100";
					when "101111100100011" => rgb <= "100100";
					when "101111100100100" => rgb <= "100100";
					when "101111100100101" => rgb <= "100100";
					when "101111100100110" => rgb <= "100100";
					when "101111100100111" => rgb <= "100100";
					when "101111100101000" => rgb <= "100100";
					when "101111100101001" => rgb <= "100100";
					when "101111100101010" => rgb <= "100100";
					when "101111100101011" => rgb <= "100100";
					when "101111100101100" => rgb <= "100100";
					when "101111100101101" => rgb <= "100100";
					when "101111100101110" => rgb <= "100100";
					when "101111100101111" => rgb <= "100100";
					when "101111100110000" => rgb <= "100100";
					when "101111100110001" => rgb <= "100100";
					when "101111100110010" => rgb <= "010000";
					when "101111100110011" => rgb <= "010000";
					when "101111100110100" => rgb <= "000000";
					when "101111100110101" => rgb <= "000000";
					when "101111100110110" => rgb <= "101111";
					when "101111100110111" => rgb <= "101111";
					when "101111100111000" => rgb <= "101111";
					when "101111100111001" => rgb <= "101111";
					when "101111100111010" => rgb <= "101111";
					when "101111100111011" => rgb <= "101111";
					when "101111100111100" => rgb <= "101111";
					when "101111100111101" => rgb <= "101111";
					when "101111100111110" => rgb <= "101111";
					when "101111100111111" => rgb <= "101111";
					when "101111101000000" => rgb <= "101111";
					when "101111101000001" => rgb <= "101111";
					when "101111101000010" => rgb <= "101111";
					when "101111101000011" => rgb <= "101111";
					when "101111101000100" => rgb <= "101111";
					when "101111101000101" => rgb <= "101111";
					when "101111101000110" => rgb <= "101111";
					when "101111101000111" => rgb <= "101111";
					when "101111101001000" => rgb <= "101111";
					when "101111101001001" => rgb <= "101111";
					when "101111101001010" => rgb <= "101111";
					when "101111101001011" => rgb <= "101111";
					when "101111101001100" => rgb <= "101111";
					when "101111101001101" => rgb <= "101111";
					when "101111101001110" => rgb <= "101111";
					when "101111101001111" => rgb <= "101111";
					when "101111101010000" => rgb <= "101111";
					when "101111101010001" => rgb <= "101111";
					when "101111101010010" => rgb <= "101111";
					when "101111101010011" => rgb <= "101111";
					when "101111101010100" => rgb <= "101111";
					when "101111101010101" => rgb <= "101111";
					when "101111101010110" => rgb <= "101111";
					when "101111101010111" => rgb <= "101111";
					when "101111101011000" => rgb <= "101111";
					when "101111101011001" => rgb <= "101111";
					when "101111101011010" => rgb <= "101111";
					when "101111101011011" => rgb <= "101111";
					when "101111101011100" => rgb <= "101111";
					when "101111101011101" => rgb <= "101111";
					when "101111101011110" => rgb <= "101111";
					when "101111101011111" => rgb <= "101111";
					when "101111101100000" => rgb <= "101111";
					when "101111101100001" => rgb <= "101111";
					when "101111101100010" => rgb <= "101111";
					when "101111101100011" => rgb <= "101111";
					when "101111101100100" => rgb <= "101111";
					when "101111101100101" => rgb <= "101111";
					when "101111101100110" => rgb <= "101111";
					when "101111101100111" => rgb <= "101111";
					when "101111101101000" => rgb <= "101111";
					when "101111101101001" => rgb <= "101111";
					when "101111101101010" => rgb <= "101111";
					when "101111101101011" => rgb <= "101111";
					when "101111101101100" => rgb <= "101111";
					when "101111101101101" => rgb <= "101111";
					when "101111101101110" => rgb <= "101111";
					when "101111101101111" => rgb <= "101111";
					when "101111101110000" => rgb <= "101111";
					when "101111101110001" => rgb <= "101111";
					when "101111101110010" => rgb <= "101111";
					when "101111101110011" => rgb <= "101111";
					when "101111101110100" => rgb <= "101111";
					when "101111101110101" => rgb <= "101111";
					when "101111101110110" => rgb <= "101111";
					when "101111101110111" => rgb <= "101111";
					when "101111101111000" => rgb <= "101111";
					when "101111101111001" => rgb <= "101111";
					when "101111101111010" => rgb <= "101111";
					when "101111101111011" => rgb <= "101111";
					when "101111101111100" => rgb <= "101111";
					when "101111101111101" => rgb <= "101111";
					when "101111101111110" => rgb <= "101111";
					when "101111101111111" => rgb <= "101111";
					when "101111110000000" => rgb <= "101111";
					when "101111110000001" => rgb <= "101111";
					when "101111110000010" => rgb <= "101111";
					when "101111110000011" => rgb <= "101111";
					when "101111110000100" => rgb <= "101111";
					when "101111110000101" => rgb <= "101111";
					when "101111110000110" => rgb <= "101111";
					when "101111110000111" => rgb <= "101111";
					when "101111110001000" => rgb <= "101111";
					when "101111110001001" => rgb <= "101111";
					when "101111110001010" => rgb <= "101111";
					when "101111110001011" => rgb <= "101111";
					when "101111110001100" => rgb <= "101111";
					when "101111110001101" => rgb <= "101111";
					when "101111110001110" => rgb <= "101111";
					when "101111110001111" => rgb <= "101111";
					when "101111110010000" => rgb <= "101111";
					when "101111110010001" => rgb <= "101111";
					when "101111110010010" => rgb <= "101111";
					when "101111110010011" => rgb <= "101111";
					when "101111110010100" => rgb <= "101111";
					when "101111110010101" => rgb <= "101111";
					when "101111110010110" => rgb <= "101111";
					when "101111110010111" => rgb <= "101111";
					when "101111110011000" => rgb <= "101111";
					when "101111110011001" => rgb <= "101111";
					when "101111110011010" => rgb <= "101111";
					when "101111110011011" => rgb <= "101111";
					when "101111110011100" => rgb <= "101111";
					when "101111110011101" => rgb <= "101111";
					when "101111110011110" => rgb <= "101111";
					when "101111110011111" => rgb <= "101111";
					when "110000000000000" => rgb <= "101111";
					when "110000000000001" => rgb <= "101111";
					when "110000000000010" => rgb <= "101111";
					when "110000000000011" => rgb <= "101111";
					when "110000000000100" => rgb <= "101111";
					when "110000000000101" => rgb <= "101111";
					when "110000000000110" => rgb <= "101111";
					when "110000000000111" => rgb <= "101111";
					when "110000000001000" => rgb <= "000010";
					when "110000000001001" => rgb <= "000010";
					when "110000000001010" => rgb <= "000010";
					when "110000000001011" => rgb <= "000010";
					when "110000000001100" => rgb <= "000010";
					when "110000000001101" => rgb <= "000010";
					when "110000000001110" => rgb <= "000010";
					when "110000000001111" => rgb <= "000010";
					when "110000000010000" => rgb <= "000010";
					when "110000000010001" => rgb <= "000010";
					when "110000000010010" => rgb <= "000010";
					when "110000000010011" => rgb <= "000010";
					when "110000000010100" => rgb <= "000010";
					when "110000000010101" => rgb <= "000010";
					when "110000000010110" => rgb <= "000010";
					when "110000000010111" => rgb <= "000010";
					when "110000000011000" => rgb <= "000010";
					when "110000000011001" => rgb <= "000010";
					when "110000000011010" => rgb <= "000010";
					when "110000000011011" => rgb <= "000010";
					when "110000000011100" => rgb <= "000010";
					when "110000000011101" => rgb <= "000010";
					when "110000000011110" => rgb <= "000010";
					when "110000000011111" => rgb <= "000010";
					when "110000000100000" => rgb <= "000010";
					when "110000000100001" => rgb <= "000010";
					when "110000000100010" => rgb <= "000010";
					when "110000000100011" => rgb <= "000010";
					when "110000000100100" => rgb <= "000010";
					when "110000000100101" => rgb <= "000010";
					when "110000000100110" => rgb <= "000010";
					when "110000000100111" => rgb <= "000010";
					when "110000000101000" => rgb <= "000010";
					when "110000000101001" => rgb <= "000010";
					when "110000000101010" => rgb <= "000010";
					when "110000000101011" => rgb <= "000010";
					when "110000000101100" => rgb <= "000010";
					when "110000000101101" => rgb <= "000010";
					when "110000000101110" => rgb <= "100100";
					when "110000000101111" => rgb <= "100100";
					when "110000000110000" => rgb <= "100100";
					when "110000000110001" => rgb <= "100100";
					when "110000000110010" => rgb <= "010000";
					when "110000000110011" => rgb <= "010000";
					when "110000000110100" => rgb <= "000000";
					when "110000000110101" => rgb <= "000000";
					when "110000000110110" => rgb <= "101111";
					when "110000000110111" => rgb <= "101111";
					when "110000000111000" => rgb <= "101111";
					when "110000000111001" => rgb <= "101111";
					when "110000000111010" => rgb <= "101111";
					when "110000000111011" => rgb <= "101111";
					when "110000000111100" => rgb <= "101111";
					when "110000000111101" => rgb <= "101111";
					when "110000000111110" => rgb <= "101111";
					when "110000000111111" => rgb <= "101111";
					when "110000001000000" => rgb <= "101111";
					when "110000001000001" => rgb <= "101111";
					when "110000001000010" => rgb <= "101111";
					when "110000001000011" => rgb <= "101111";
					when "110000001000100" => rgb <= "101111";
					when "110000001000101" => rgb <= "101111";
					when "110000001000110" => rgb <= "101111";
					when "110000001000111" => rgb <= "101111";
					when "110000001001000" => rgb <= "101111";
					when "110000001001001" => rgb <= "101111";
					when "110000001001010" => rgb <= "101111";
					when "110000001001011" => rgb <= "101111";
					when "110000001001100" => rgb <= "101111";
					when "110000001001101" => rgb <= "101111";
					when "110000001001110" => rgb <= "101111";
					when "110000001001111" => rgb <= "101111";
					when "110000001010000" => rgb <= "101111";
					when "110000001010001" => rgb <= "101111";
					when "110000001010010" => rgb <= "101111";
					when "110000001010011" => rgb <= "101111";
					when "110000001010100" => rgb <= "101111";
					when "110000001010101" => rgb <= "101111";
					when "110000001010110" => rgb <= "101111";
					when "110000001010111" => rgb <= "101111";
					when "110000001011000" => rgb <= "101111";
					when "110000001011001" => rgb <= "101111";
					when "110000001011010" => rgb <= "101111";
					when "110000001011011" => rgb <= "101111";
					when "110000001011100" => rgb <= "101111";
					when "110000001011101" => rgb <= "101111";
					when "110000001011110" => rgb <= "101111";
					when "110000001011111" => rgb <= "101111";
					when "110000001100000" => rgb <= "101111";
					when "110000001100001" => rgb <= "101111";
					when "110000001100010" => rgb <= "101111";
					when "110000001100011" => rgb <= "101111";
					when "110000001100100" => rgb <= "101111";
					when "110000001100101" => rgb <= "101111";
					when "110000001100110" => rgb <= "101111";
					when "110000001100111" => rgb <= "101111";
					when "110000001101000" => rgb <= "101111";
					when "110000001101001" => rgb <= "101111";
					when "110000001101010" => rgb <= "101111";
					when "110000001101011" => rgb <= "101111";
					when "110000001101100" => rgb <= "101111";
					when "110000001101101" => rgb <= "101111";
					when "110000001101110" => rgb <= "101111";
					when "110000001101111" => rgb <= "101111";
					when "110000001110000" => rgb <= "101111";
					when "110000001110001" => rgb <= "101111";
					when "110000001110010" => rgb <= "000010";
					when "110000001110011" => rgb <= "000010";
					when "110000001110100" => rgb <= "000010";
					when "110000001110101" => rgb <= "000010";
					when "110000001110110" => rgb <= "000010";
					when "110000001110111" => rgb <= "000010";
					when "110000001111000" => rgb <= "000010";
					when "110000001111001" => rgb <= "000010";
					when "110000001111010" => rgb <= "000010";
					when "110000001111011" => rgb <= "000010";
					when "110000001111100" => rgb <= "000010";
					when "110000001111101" => rgb <= "000010";
					when "110000001111110" => rgb <= "000010";
					when "110000001111111" => rgb <= "000010";
					when "110000010000000" => rgb <= "000010";
					when "110000010000001" => rgb <= "000010";
					when "110000010000010" => rgb <= "000010";
					when "110000010000011" => rgb <= "000010";
					when "110000010000100" => rgb <= "000010";
					when "110000010000101" => rgb <= "000010";
					when "110000010000110" => rgb <= "000010";
					when "110000010000111" => rgb <= "000010";
					when "110000010001000" => rgb <= "000010";
					when "110000010001001" => rgb <= "000010";
					when "110000010001010" => rgb <= "000010";
					when "110000010001011" => rgb <= "000010";
					when "110000010001100" => rgb <= "000010";
					when "110000010001101" => rgb <= "000010";
					when "110000010001110" => rgb <= "000010";
					when "110000010001111" => rgb <= "000010";
					when "110000010010000" => rgb <= "000010";
					when "110000010010001" => rgb <= "000010";
					when "110000010010010" => rgb <= "000010";
					when "110000010010011" => rgb <= "000010";
					when "110000010010100" => rgb <= "000010";
					when "110000010010101" => rgb <= "000010";
					when "110000010010110" => rgb <= "000010";
					when "110000010010111" => rgb <= "000010";
					when "110000010011000" => rgb <= "101111";
					when "110000010011001" => rgb <= "101111";
					when "110000010011010" => rgb <= "101111";
					when "110000010011011" => rgb <= "101111";
					when "110000010011100" => rgb <= "101111";
					when "110000010011101" => rgb <= "101111";
					when "110000010011110" => rgb <= "101111";
					when "110000010011111" => rgb <= "101111";
					when "110000100000000" => rgb <= "101111";
					when "110000100000001" => rgb <= "101111";
					when "110000100000010" => rgb <= "101111";
					when "110000100000011" => rgb <= "101111";
					when "110000100000100" => rgb <= "101111";
					when "110000100000101" => rgb <= "101111";
					when "110000100000110" => rgb <= "101111";
					when "110000100000111" => rgb <= "101111";
					when "110000100001000" => rgb <= "000010";
					when "110000100001001" => rgb <= "000010";
					when "110000100001010" => rgb <= "000010";
					when "110000100001011" => rgb <= "000010";
					when "110000100001100" => rgb <= "000010";
					when "110000100001101" => rgb <= "000010";
					when "110000100001110" => rgb <= "000010";
					when "110000100001111" => rgb <= "000010";
					when "110000100010000" => rgb <= "000010";
					when "110000100010001" => rgb <= "000010";
					when "110000100010010" => rgb <= "000010";
					when "110000100010011" => rgb <= "000010";
					when "110000100010100" => rgb <= "000010";
					when "110000100010101" => rgb <= "000010";
					when "110000100010110" => rgb <= "000010";
					when "110000100010111" => rgb <= "000010";
					when "110000100011000" => rgb <= "000010";
					when "110000100011001" => rgb <= "000010";
					when "110000100011010" => rgb <= "000010";
					when "110000100011011" => rgb <= "000010";
					when "110000100011100" => rgb <= "000010";
					when "110000100011101" => rgb <= "000010";
					when "110000100011110" => rgb <= "000010";
					when "110000100011111" => rgb <= "000010";
					when "110000100100000" => rgb <= "000010";
					when "110000100100001" => rgb <= "000010";
					when "110000100100010" => rgb <= "000010";
					when "110000100100011" => rgb <= "000010";
					when "110000100100100" => rgb <= "000010";
					when "110000100100101" => rgb <= "000010";
					when "110000100100110" => rgb <= "000010";
					when "110000100100111" => rgb <= "000010";
					when "110000100101000" => rgb <= "000010";
					when "110000100101001" => rgb <= "000010";
					when "110000100101010" => rgb <= "000010";
					when "110000100101011" => rgb <= "000010";
					when "110000100101100" => rgb <= "000010";
					when "110000100101101" => rgb <= "000010";
					when "110000100101110" => rgb <= "100100";
					when "110000100101111" => rgb <= "100100";
					when "110000100110000" => rgb <= "100100";
					when "110000100110001" => rgb <= "100100";
					when "110000100110010" => rgb <= "010000";
					when "110000100110011" => rgb <= "010000";
					when "110000100110100" => rgb <= "000000";
					when "110000100110101" => rgb <= "000000";
					when "110000100110110" => rgb <= "101111";
					when "110000100110111" => rgb <= "101111";
					when "110000100111000" => rgb <= "101111";
					when "110000100111001" => rgb <= "101111";
					when "110000100111010" => rgb <= "101111";
					when "110000100111011" => rgb <= "101111";
					when "110000100111100" => rgb <= "101111";
					when "110000100111101" => rgb <= "101111";
					when "110000100111110" => rgb <= "101111";
					when "110000100111111" => rgb <= "101111";
					when "110000101000000" => rgb <= "101111";
					when "110000101000001" => rgb <= "101111";
					when "110000101000010" => rgb <= "101111";
					when "110000101000011" => rgb <= "101111";
					when "110000101000100" => rgb <= "101111";
					when "110000101000101" => rgb <= "101111";
					when "110000101000110" => rgb <= "101111";
					when "110000101000111" => rgb <= "101111";
					when "110000101001000" => rgb <= "101111";
					when "110000101001001" => rgb <= "101111";
					when "110000101001010" => rgb <= "101111";
					when "110000101001011" => rgb <= "101111";
					when "110000101001100" => rgb <= "101111";
					when "110000101001101" => rgb <= "101111";
					when "110000101001110" => rgb <= "101111";
					when "110000101001111" => rgb <= "101111";
					when "110000101010000" => rgb <= "101111";
					when "110000101010001" => rgb <= "101111";
					when "110000101010010" => rgb <= "101111";
					when "110000101010011" => rgb <= "101111";
					when "110000101010100" => rgb <= "101111";
					when "110000101010101" => rgb <= "101111";
					when "110000101010110" => rgb <= "101111";
					when "110000101010111" => rgb <= "101111";
					when "110000101011000" => rgb <= "101111";
					when "110000101011001" => rgb <= "101111";
					when "110000101011010" => rgb <= "101111";
					when "110000101011011" => rgb <= "101111";
					when "110000101011100" => rgb <= "101111";
					when "110000101011101" => rgb <= "101111";
					when "110000101011110" => rgb <= "101111";
					when "110000101011111" => rgb <= "101111";
					when "110000101100000" => rgb <= "101111";
					when "110000101100001" => rgb <= "101111";
					when "110000101100010" => rgb <= "101111";
					when "110000101100011" => rgb <= "101111";
					when "110000101100100" => rgb <= "101111";
					when "110000101100101" => rgb <= "101111";
					when "110000101100110" => rgb <= "101111";
					when "110000101100111" => rgb <= "101111";
					when "110000101101000" => rgb <= "101111";
					when "110000101101001" => rgb <= "101111";
					when "110000101101010" => rgb <= "101111";
					when "110000101101011" => rgb <= "101111";
					when "110000101101100" => rgb <= "101111";
					when "110000101101101" => rgb <= "101111";
					when "110000101101110" => rgb <= "101111";
					when "110000101101111" => rgb <= "101111";
					when "110000101110000" => rgb <= "101111";
					when "110000101110001" => rgb <= "101111";
					when "110000101110010" => rgb <= "000010";
					when "110000101110011" => rgb <= "000010";
					when "110000101110100" => rgb <= "000010";
					when "110000101110101" => rgb <= "000010";
					when "110000101110110" => rgb <= "000010";
					when "110000101110111" => rgb <= "000010";
					when "110000101111000" => rgb <= "000010";
					when "110000101111001" => rgb <= "000010";
					when "110000101111010" => rgb <= "000010";
					when "110000101111011" => rgb <= "000010";
					when "110000101111100" => rgb <= "000010";
					when "110000101111101" => rgb <= "000010";
					when "110000101111110" => rgb <= "000010";
					when "110000101111111" => rgb <= "000010";
					when "110000110000000" => rgb <= "000010";
					when "110000110000001" => rgb <= "000010";
					when "110000110000010" => rgb <= "000010";
					when "110000110000011" => rgb <= "000010";
					when "110000110000100" => rgb <= "000010";
					when "110000110000101" => rgb <= "000010";
					when "110000110000110" => rgb <= "000010";
					when "110000110000111" => rgb <= "000010";
					when "110000110001000" => rgb <= "000010";
					when "110000110001001" => rgb <= "000010";
					when "110000110001010" => rgb <= "000010";
					when "110000110001011" => rgb <= "000010";
					when "110000110001100" => rgb <= "000010";
					when "110000110001101" => rgb <= "000010";
					when "110000110001110" => rgb <= "000010";
					when "110000110001111" => rgb <= "000010";
					when "110000110010000" => rgb <= "000010";
					when "110000110010001" => rgb <= "000010";
					when "110000110010010" => rgb <= "000010";
					when "110000110010011" => rgb <= "000010";
					when "110000110010100" => rgb <= "000010";
					when "110000110010101" => rgb <= "000010";
					when "110000110010110" => rgb <= "000010";
					when "110000110010111" => rgb <= "000010";
					when "110000110011000" => rgb <= "101111";
					when "110000110011001" => rgb <= "101111";
					when "110000110011010" => rgb <= "101111";
					when "110000110011011" => rgb <= "101111";
					when "110000110011100" => rgb <= "101111";
					when "110000110011101" => rgb <= "101111";
					when "110000110011110" => rgb <= "101111";
					when "110000110011111" => rgb <= "101111";
					when "110001000000000" => rgb <= "101111";
					when "110001000000001" => rgb <= "101111";
					when "110001000000010" => rgb <= "101111";
					when "110001000000011" => rgb <= "101111";
					when "110001000000100" => rgb <= "101111";
					when "110001000000101" => rgb <= "101111";
					when "110001000000110" => rgb <= "101111";
					when "110001000000111" => rgb <= "101111";
					when "110001000001000" => rgb <= "000011";
					when "110001000001001" => rgb <= "000011";
					when "110001000001010" => rgb <= "000011";
					when "110001000001011" => rgb <= "000011";
					when "110001000001100" => rgb <= "000011";
					when "110001000001101" => rgb <= "000011";
					when "110001000001110" => rgb <= "000011";
					when "110001000001111" => rgb <= "000011";
					when "110001000010000" => rgb <= "000011";
					when "110001000010001" => rgb <= "000011";
					when "110001000010010" => rgb <= "000011";
					when "110001000010011" => rgb <= "000011";
					when "110001000010100" => rgb <= "000011";
					when "110001000010101" => rgb <= "000011";
					when "110001000010110" => rgb <= "000011";
					when "110001000010111" => rgb <= "101111";
					when "110001000011000" => rgb <= "000011";
					when "110001000011001" => rgb <= "000011";
					when "110001000011010" => rgb <= "000011";
					when "110001000011011" => rgb <= "000011";
					when "110001000011100" => rgb <= "000011";
					when "110001000011101" => rgb <= "000011";
					when "110001000011110" => rgb <= "000011";
					when "110001000011111" => rgb <= "000011";
					when "110001000100000" => rgb <= "000011";
					when "110001000100001" => rgb <= "000011";
					when "110001000100010" => rgb <= "000011";
					when "110001000100011" => rgb <= "000011";
					when "110001000100100" => rgb <= "000011";
					when "110001000100101" => rgb <= "000011";
					when "110001000100110" => rgb <= "000011";
					when "110001000100111" => rgb <= "000011";
					when "110001000101000" => rgb <= "000011";
					when "110001000101001" => rgb <= "000011";
					when "110001000101010" => rgb <= "000011";
					when "110001000101011" => rgb <= "000011";
					when "110001000101100" => rgb <= "000011";
					when "110001000101101" => rgb <= "000011";
					when "110001000101110" => rgb <= "100100";
					when "110001000101111" => rgb <= "100100";
					when "110001000110000" => rgb <= "100100";
					when "110001000110001" => rgb <= "100100";
					when "110001000110010" => rgb <= "010000";
					when "110001000110011" => rgb <= "010000";
					when "110001000110100" => rgb <= "000000";
					when "110001000110101" => rgb <= "000000";
					when "110001000110110" => rgb <= "101111";
					when "110001000110111" => rgb <= "101111";
					when "110001000111000" => rgb <= "101111";
					when "110001000111001" => rgb <= "101111";
					when "110001000111010" => rgb <= "101111";
					when "110001000111011" => rgb <= "101111";
					when "110001000111100" => rgb <= "101111";
					when "110001000111101" => rgb <= "101111";
					when "110001000111110" => rgb <= "101111";
					when "110001000111111" => rgb <= "101111";
					when "110001001000000" => rgb <= "101111";
					when "110001001000001" => rgb <= "101111";
					when "110001001000010" => rgb <= "101111";
					when "110001001000011" => rgb <= "101111";
					when "110001001000100" => rgb <= "101111";
					when "110001001000101" => rgb <= "101111";
					when "110001001000110" => rgb <= "101111";
					when "110001001000111" => rgb <= "101111";
					when "110001001001000" => rgb <= "101111";
					when "110001001001001" => rgb <= "101111";
					when "110001001001010" => rgb <= "101111";
					when "110001001001011" => rgb <= "101111";
					when "110001001001100" => rgb <= "101111";
					when "110001001001101" => rgb <= "101111";
					when "110001001001110" => rgb <= "101111";
					when "110001001001111" => rgb <= "101111";
					when "110001001010000" => rgb <= "101111";
					when "110001001010001" => rgb <= "101111";
					when "110001001010010" => rgb <= "101111";
					when "110001001010011" => rgb <= "101111";
					when "110001001010100" => rgb <= "101111";
					when "110001001010101" => rgb <= "101111";
					when "110001001010110" => rgb <= "101111";
					when "110001001010111" => rgb <= "101111";
					when "110001001011000" => rgb <= "101111";
					when "110001001011001" => rgb <= "101111";
					when "110001001011010" => rgb <= "101111";
					when "110001001011011" => rgb <= "101111";
					when "110001001011100" => rgb <= "101111";
					when "110001001011101" => rgb <= "101111";
					when "110001001011110" => rgb <= "101111";
					when "110001001011111" => rgb <= "101111";
					when "110001001100000" => rgb <= "101111";
					when "110001001100001" => rgb <= "101111";
					when "110001001100010" => rgb <= "101111";
					when "110001001100011" => rgb <= "101111";
					when "110001001100100" => rgb <= "101111";
					when "110001001100101" => rgb <= "101111";
					when "110001001100110" => rgb <= "101111";
					when "110001001100111" => rgb <= "101111";
					when "110001001101000" => rgb <= "101111";
					when "110001001101001" => rgb <= "101111";
					when "110001001101010" => rgb <= "101111";
					when "110001001101011" => rgb <= "101111";
					when "110001001101100" => rgb <= "101111";
					when "110001001101101" => rgb <= "101111";
					when "110001001101110" => rgb <= "101111";
					when "110001001101111" => rgb <= "101111";
					when "110001001110000" => rgb <= "101111";
					when "110001001110001" => rgb <= "101111";
					when "110001001110010" => rgb <= "000011";
					when "110001001110011" => rgb <= "000011";
					when "110001001110100" => rgb <= "000011";
					when "110001001110101" => rgb <= "000011";
					when "110001001110110" => rgb <= "000011";
					when "110001001110111" => rgb <= "000011";
					when "110001001111000" => rgb <= "101111";
					when "110001001111001" => rgb <= "101111";
					when "110001001111010" => rgb <= "000011";
					when "110001001111011" => rgb <= "000011";
					when "110001001111100" => rgb <= "000011";
					when "110001001111101" => rgb <= "000011";
					when "110001001111110" => rgb <= "000011";
					when "110001001111111" => rgb <= "000011";
					when "110001010000000" => rgb <= "000011";
					when "110001010000001" => rgb <= "000011";
					when "110001010000010" => rgb <= "000011";
					when "110001010000011" => rgb <= "000011";
					when "110001010000100" => rgb <= "000011";
					when "110001010000101" => rgb <= "000011";
					when "110001010000110" => rgb <= "000011";
					when "110001010000111" => rgb <= "000011";
					when "110001010001000" => rgb <= "000011";
					when "110001010001001" => rgb <= "000011";
					when "110001010001010" => rgb <= "000011";
					when "110001010001011" => rgb <= "000011";
					when "110001010001100" => rgb <= "000011";
					when "110001010001101" => rgb <= "000011";
					when "110001010001110" => rgb <= "000011";
					when "110001010001111" => rgb <= "000011";
					when "110001010010000" => rgb <= "000011";
					when "110001010010001" => rgb <= "000011";
					when "110001010010010" => rgb <= "000011";
					when "110001010010011" => rgb <= "000011";
					when "110001010010100" => rgb <= "000011";
					when "110001010010101" => rgb <= "000011";
					when "110001010010110" => rgb <= "000011";
					when "110001010010111" => rgb <= "000011";
					when "110001010011000" => rgb <= "101111";
					when "110001010011001" => rgb <= "101111";
					when "110001010011010" => rgb <= "101111";
					when "110001010011011" => rgb <= "101111";
					when "110001010011100" => rgb <= "101111";
					when "110001010011101" => rgb <= "101111";
					when "110001010011110" => rgb <= "101111";
					when "110001010011111" => rgb <= "101111";
					when "110001100000000" => rgb <= "101111";
					when "110001100000001" => rgb <= "101111";
					when "110001100000010" => rgb <= "101111";
					when "110001100000011" => rgb <= "101111";
					when "110001100000100" => rgb <= "101111";
					when "110001100000101" => rgb <= "101111";
					when "110001100000110" => rgb <= "101111";
					when "110001100000111" => rgb <= "101111";
					when "110001100001000" => rgb <= "101111";
					when "110001100001001" => rgb <= "000011";
					when "110001100001010" => rgb <= "000011";
					when "110001100001011" => rgb <= "101111";
					when "110001100001100" => rgb <= "000011";
					when "110001100001101" => rgb <= "101111";
					when "110001100001110" => rgb <= "101111";
					when "110001100001111" => rgb <= "101111";
					when "110001100010000" => rgb <= "000011";
					when "110001100010001" => rgb <= "101111";
					when "110001100010010" => rgb <= "000011";
					when "110001100010011" => rgb <= "000011";
					when "110001100010100" => rgb <= "101111";
					when "110001100010101" => rgb <= "000011";
					when "110001100010110" => rgb <= "101111";
					when "110001100010111" => rgb <= "101111";
					when "110001100011000" => rgb <= "101111";
					when "110001100011001" => rgb <= "000011";
					when "110001100011010" => rgb <= "000011";
					when "110001100011011" => rgb <= "000011";
					when "110001100011100" => rgb <= "101111";
					when "110001100011101" => rgb <= "101111";
					when "110001100011110" => rgb <= "000011";
					when "110001100011111" => rgb <= "101111";
					when "110001100100000" => rgb <= "000000";
					when "110001100100001" => rgb <= "000011";
					when "110001100100010" => rgb <= "100100";
					when "110001100100011" => rgb <= "100100";
					when "110001100100100" => rgb <= "100100";
					when "110001100100101" => rgb <= "000011";
					when "110001100100110" => rgb <= "100100";
					when "110001100100111" => rgb <= "000011";
					when "110001100101000" => rgb <= "100100";
					when "110001100101001" => rgb <= "000011";
					when "110001100101010" => rgb <= "000011";
					when "110001100101011" => rgb <= "000011";
					when "110001100101100" => rgb <= "000011";
					when "110001100101101" => rgb <= "100100";
					when "110001100101110" => rgb <= "100100";
					when "110001100101111" => rgb <= "100100";
					when "110001100110000" => rgb <= "100100";
					when "110001100110001" => rgb <= "100100";
					when "110001100110010" => rgb <= "010000";
					when "110001100110011" => rgb <= "010000";
					when "110001100110100" => rgb <= "000000";
					when "110001100110101" => rgb <= "000000";
					when "110001100110110" => rgb <= "101111";
					when "110001100110111" => rgb <= "101111";
					when "110001100111000" => rgb <= "101111";
					when "110001100111001" => rgb <= "101111";
					when "110001100111010" => rgb <= "101111";
					when "110001100111011" => rgb <= "101111";
					when "110001100111100" => rgb <= "101111";
					when "110001100111101" => rgb <= "101111";
					when "110001100111110" => rgb <= "101111";
					when "110001100111111" => rgb <= "101111";
					when "110001101000000" => rgb <= "101111";
					when "110001101000001" => rgb <= "101111";
					when "110001101000010" => rgb <= "101111";
					when "110001101000011" => rgb <= "101111";
					when "110001101000100" => rgb <= "101111";
					when "110001101000101" => rgb <= "101111";
					when "110001101000110" => rgb <= "101111";
					when "110001101000111" => rgb <= "101111";
					when "110001101001000" => rgb <= "101111";
					when "110001101001001" => rgb <= "101111";
					when "110001101001010" => rgb <= "101111";
					when "110001101001011" => rgb <= "101111";
					when "110001101001100" => rgb <= "101111";
					when "110001101001101" => rgb <= "101111";
					when "110001101001110" => rgb <= "101111";
					when "110001101001111" => rgb <= "101111";
					when "110001101010000" => rgb <= "101111";
					when "110001101010001" => rgb <= "101111";
					when "110001101010010" => rgb <= "101111";
					when "110001101010011" => rgb <= "101111";
					when "110001101010100" => rgb <= "101111";
					when "110001101010101" => rgb <= "101111";
					when "110001101010110" => rgb <= "101111";
					when "110001101010111" => rgb <= "101111";
					when "110001101011000" => rgb <= "101111";
					when "110001101011001" => rgb <= "101111";
					when "110001101011010" => rgb <= "101111";
					when "110001101011011" => rgb <= "101111";
					when "110001101011100" => rgb <= "101111";
					when "110001101011101" => rgb <= "101111";
					when "110001101011110" => rgb <= "101111";
					when "110001101011111" => rgb <= "101111";
					when "110001101100000" => rgb <= "101111";
					when "110001101100001" => rgb <= "101111";
					when "110001101100010" => rgb <= "101111";
					when "110001101100011" => rgb <= "101111";
					when "110001101100100" => rgb <= "101111";
					when "110001101100101" => rgb <= "101111";
					when "110001101100110" => rgb <= "101111";
					when "110001101100111" => rgb <= "101111";
					when "110001101101000" => rgb <= "101111";
					when "110001101101001" => rgb <= "101111";
					when "110001101101010" => rgb <= "101111";
					when "110001101101011" => rgb <= "101111";
					when "110001101101100" => rgb <= "101111";
					when "110001101101101" => rgb <= "101111";
					when "110001101101110" => rgb <= "101111";
					when "110001101101111" => rgb <= "101111";
					when "110001101110000" => rgb <= "101111";
					when "110001101110001" => rgb <= "101111";
					when "110001101110010" => rgb <= "101111";
					when "110001101110011" => rgb <= "000011";
					when "110001101110100" => rgb <= "000011";
					when "110001101110101" => rgb <= "000011";
					when "110001101110110" => rgb <= "101111";
					when "110001101110111" => rgb <= "101111";
					when "110001101111000" => rgb <= "101111";
					when "110001101111001" => rgb <= "101111";
					when "110001101111010" => rgb <= "101111";
					when "110001101111011" => rgb <= "101111";
					when "110001101111100" => rgb <= "000011";
					when "110001101111101" => rgb <= "000011";
					when "110001101111110" => rgb <= "000011";
					when "110001101111111" => rgb <= "000011";
					when "110001110000000" => rgb <= "000011";
					when "110001110000001" => rgb <= "000011";
					when "110001110000010" => rgb <= "101111";
					when "110001110000011" => rgb <= "000011";
					when "110001110000100" => rgb <= "000011";
					when "110001110000101" => rgb <= "000011";
					when "110001110000110" => rgb <= "101111";
					when "110001110000111" => rgb <= "101111";
					when "110001110001000" => rgb <= "000011";
					when "110001110001001" => rgb <= "000011";
					when "110001110001010" => rgb <= "000011";
					when "110001110001011" => rgb <= "000011";
					when "110001110001100" => rgb <= "000011";
					when "110001110001101" => rgb <= "000011";
					when "110001110001110" => rgb <= "000011";
					when "110001110001111" => rgb <= "101111";
					when "110001110010000" => rgb <= "101111";
					when "110001110010001" => rgb <= "000011";
					when "110001110010010" => rgb <= "000011";
					when "110001110010011" => rgb <= "101111";
					when "110001110010100" => rgb <= "000011";
					when "110001110010101" => rgb <= "000011";
					when "110001110010110" => rgb <= "101111";
					when "110001110010111" => rgb <= "101111";
					when "110001110011000" => rgb <= "101111";
					when "110001110011001" => rgb <= "101111";
					when "110001110011010" => rgb <= "101111";
					when "110001110011011" => rgb <= "101111";
					when "110001110011100" => rgb <= "101111";
					when "110001110011101" => rgb <= "101111";
					when "110001110011110" => rgb <= "101111";
					when "110001110011111" => rgb <= "101111";
					when "110010000000000" => rgb <= "101111";
					when "110010000000001" => rgb <= "101111";
					when "110010000000010" => rgb <= "101111";
					when "110010000000011" => rgb <= "101111";
					when "110010000000100" => rgb <= "101111";
					when "110010000000101" => rgb <= "101111";
					when "110010000000110" => rgb <= "101111";
					when "110010000000111" => rgb <= "101111";
					when "110010000001000" => rgb <= "101111";
					when "110010000001001" => rgb <= "101111";
					when "110010000001010" => rgb <= "000011";
					when "110010000001011" => rgb <= "101111";
					when "110010000001100" => rgb <= "101111";
					when "110010000001101" => rgb <= "101111";
					when "110010000001110" => rgb <= "101111";
					when "110010000001111" => rgb <= "101111";
					when "110010000010000" => rgb <= "101111";
					when "110010000010001" => rgb <= "101111";
					when "110010000010010" => rgb <= "000011";
					when "110010000010011" => rgb <= "101111";
					when "110010000010100" => rgb <= "101111";
					when "110010000010101" => rgb <= "101111";
					when "110010000010110" => rgb <= "101111";
					when "110010000010111" => rgb <= "101111";
					when "110010000011000" => rgb <= "101111";
					when "110010000011001" => rgb <= "101111";
					when "110010000011010" => rgb <= "101111";
					when "110010000011011" => rgb <= "000011";
					when "110010000011100" => rgb <= "101111";
					when "110010000011101" => rgb <= "101111";
					when "110010000011110" => rgb <= "000000";
					when "110010000011111" => rgb <= "000000";
					when "110010000100000" => rgb <= "100100";
					when "110010000100001" => rgb <= "100100";
					when "110010000100010" => rgb <= "100100";
					when "110010000100011" => rgb <= "100100";
					when "110010000100100" => rgb <= "100100";
					when "110010000100101" => rgb <= "100100";
					when "110010000100110" => rgb <= "100100";
					when "110010000100111" => rgb <= "100100";
					when "110010000101000" => rgb <= "100100";
					when "110010000101001" => rgb <= "000011";
					when "110010000101010" => rgb <= "000011";
					when "110010000101011" => rgb <= "000011";
					when "110010000101100" => rgb <= "100100";
					when "110010000101101" => rgb <= "100100";
					when "110010000101110" => rgb <= "100100";
					when "110010000101111" => rgb <= "100100";
					when "110010000110000" => rgb <= "100100";
					when "110010000110001" => rgb <= "100100";
					when "110010000110010" => rgb <= "010000";
					when "110010000110011" => rgb <= "010000";
					when "110010000110100" => rgb <= "000000";
					when "110010000110101" => rgb <= "000000";
					when "110010000110110" => rgb <= "000000";
					when "110010000110111" => rgb <= "000000";
					when "110010000111000" => rgb <= "101111";
					when "110010000111001" => rgb <= "101111";
					when "110010000111010" => rgb <= "101111";
					when "110010000111011" => rgb <= "101111";
					when "110010000111100" => rgb <= "101111";
					when "110010000111101" => rgb <= "101111";
					when "110010000111110" => rgb <= "101111";
					when "110010000111111" => rgb <= "101111";
					when "110010001000000" => rgb <= "101111";
					when "110010001000001" => rgb <= "101111";
					when "110010001000010" => rgb <= "101111";
					when "110010001000011" => rgb <= "101111";
					when "110010001000100" => rgb <= "101111";
					when "110010001000101" => rgb <= "101111";
					when "110010001000110" => rgb <= "101111";
					when "110010001000111" => rgb <= "101111";
					when "110010001001000" => rgb <= "101111";
					when "110010001001001" => rgb <= "101111";
					when "110010001001010" => rgb <= "101111";
					when "110010001001011" => rgb <= "101111";
					when "110010001001100" => rgb <= "101111";
					when "110010001001101" => rgb <= "101111";
					when "110010001001110" => rgb <= "101111";
					when "110010001001111" => rgb <= "101111";
					when "110010001010000" => rgb <= "101111";
					when "110010001010001" => rgb <= "101111";
					when "110010001010010" => rgb <= "101111";
					when "110010001010011" => rgb <= "101111";
					when "110010001010100" => rgb <= "101111";
					when "110010001010101" => rgb <= "101111";
					when "110010001010110" => rgb <= "101111";
					when "110010001010111" => rgb <= "101111";
					when "110010001011000" => rgb <= "101111";
					when "110010001011001" => rgb <= "101111";
					when "110010001011010" => rgb <= "101111";
					when "110010001011011" => rgb <= "101111";
					when "110010001011100" => rgb <= "101111";
					when "110010001011101" => rgb <= "101111";
					when "110010001011110" => rgb <= "101111";
					when "110010001011111" => rgb <= "101111";
					when "110010001100000" => rgb <= "101111";
					when "110010001100001" => rgb <= "101111";
					when "110010001100010" => rgb <= "101111";
					when "110010001100011" => rgb <= "101111";
					when "110010001100100" => rgb <= "101111";
					when "110010001100101" => rgb <= "101111";
					when "110010001100110" => rgb <= "101111";
					when "110010001100111" => rgb <= "101111";
					when "110010001101000" => rgb <= "101111";
					when "110010001101001" => rgb <= "101111";
					when "110010001101010" => rgb <= "101111";
					when "110010001101011" => rgb <= "101111";
					when "110010001101100" => rgb <= "101111";
					when "110010001101101" => rgb <= "101111";
					when "110010001101110" => rgb <= "101111";
					when "110010001101111" => rgb <= "101111";
					when "110010001110000" => rgb <= "101111";
					when "110010001110001" => rgb <= "101111";
					when "110010001110010" => rgb <= "101111";
					when "110010001110011" => rgb <= "101111";
					when "110010001110100" => rgb <= "101111";
					when "110010001110101" => rgb <= "000011";
					when "110010001110110" => rgb <= "101111";
					when "110010001110111" => rgb <= "101111";
					when "110010001111000" => rgb <= "101111";
					when "110010001111001" => rgb <= "101111";
					when "110010001111010" => rgb <= "101111";
					when "110010001111011" => rgb <= "101111";
					when "110010001111100" => rgb <= "101111";
					when "110010001111101" => rgb <= "101111";
					when "110010001111110" => rgb <= "000011";
					when "110010001111111" => rgb <= "101111";
					when "110010010000000" => rgb <= "101111";
					when "110010010000001" => rgb <= "000011";
					when "110010010000010" => rgb <= "101111";
					when "110010010000011" => rgb <= "101111";
					when "110010010000100" => rgb <= "101111";
					when "110010010000101" => rgb <= "000011";
					when "110010010000110" => rgb <= "101111";
					when "110010010000111" => rgb <= "101111";
					when "110010010001000" => rgb <= "101111";
					when "110010010001001" => rgb <= "101111";
					when "110010010001010" => rgb <= "000011";
					when "110010010001011" => rgb <= "000011";
					when "110010010001100" => rgb <= "000011";
					when "110010010001101" => rgb <= "101111";
					when "110010010001110" => rgb <= "101111";
					when "110010010001111" => rgb <= "101111";
					when "110010010010000" => rgb <= "101111";
					when "110010010010001" => rgb <= "101111";
					when "110010010010010" => rgb <= "101111";
					when "110010010010011" => rgb <= "101111";
					when "110010010010100" => rgb <= "101111";
					when "110010010010101" => rgb <= "101111";
					when "110010010010110" => rgb <= "101111";
					when "110010010010111" => rgb <= "101111";
					when "110010010011000" => rgb <= "101111";
					when "110010010011001" => rgb <= "101111";
					when "110010010011010" => rgb <= "101111";
					when "110010010011011" => rgb <= "101111";
					when "110010010011100" => rgb <= "101111";
					when "110010010011101" => rgb <= "101111";
					when "110010010011110" => rgb <= "101111";
					when "110010010011111" => rgb <= "101111";
					when "110010100000000" => rgb <= "101111";
					when "110010100000001" => rgb <= "101111";
					when "110010100000010" => rgb <= "101111";
					when "110010100000011" => rgb <= "101111";
					when "110010100000100" => rgb <= "101111";
					when "110010100000101" => rgb <= "101111";
					when "110010100000110" => rgb <= "101111";
					when "110010100000111" => rgb <= "101111";
					when "110010100001000" => rgb <= "101111";
					when "110010100001001" => rgb <= "101111";
					when "110010100001010" => rgb <= "101111";
					when "110010100001011" => rgb <= "101111";
					when "110010100001100" => rgb <= "101111";
					when "110010100001101" => rgb <= "101111";
					when "110010100001110" => rgb <= "101111";
					when "110010100001111" => rgb <= "101111";
					when "110010100010000" => rgb <= "101111";
					when "110010100010001" => rgb <= "101111";
					when "110010100010010" => rgb <= "101111";
					when "110010100010011" => rgb <= "101111";
					when "110010100010100" => rgb <= "101111";
					when "110010100010101" => rgb <= "101111";
					when "110010100010110" => rgb <= "101111";
					when "110010100010111" => rgb <= "101111";
					when "110010100011000" => rgb <= "101111";
					when "110010100011001" => rgb <= "101111";
					when "110010100011010" => rgb <= "101111";
					when "110010100011011" => rgb <= "101111";
					when "110010100011100" => rgb <= "101111";
					when "110010100011101" => rgb <= "101111";
					when "110010100011110" => rgb <= "000000";
					when "110010100011111" => rgb <= "000000";
					when "110010100100000" => rgb <= "100100";
					when "110010100100001" => rgb <= "100100";
					when "110010100100010" => rgb <= "100100";
					when "110010100100011" => rgb <= "100100";
					when "110010100100100" => rgb <= "100100";
					when "110010100100101" => rgb <= "100100";
					when "110010100100110" => rgb <= "100100";
					when "110010100100111" => rgb <= "100100";
					when "110010100101000" => rgb <= "100100";
					when "110010100101001" => rgb <= "100100";
					when "110010100101010" => rgb <= "100100";
					when "110010100101011" => rgb <= "000011";
					when "110010100101100" => rgb <= "100100";
					when "110010100101101" => rgb <= "100100";
					when "110010100101110" => rgb <= "100100";
					when "110010100101111" => rgb <= "100100";
					when "110010100110000" => rgb <= "100100";
					when "110010100110001" => rgb <= "100100";
					when "110010100110010" => rgb <= "010000";
					when "110010100110011" => rgb <= "010000";
					when "110010100110100" => rgb <= "000000";
					when "110010100110101" => rgb <= "000000";
					when "110010100110110" => rgb <= "000000";
					when "110010100110111" => rgb <= "000000";
					when "110010100111000" => rgb <= "101111";
					when "110010100111001" => rgb <= "101111";
					when "110010100111010" => rgb <= "101111";
					when "110010100111011" => rgb <= "101111";
					when "110010100111100" => rgb <= "101111";
					when "110010100111101" => rgb <= "101111";
					when "110010100111110" => rgb <= "101111";
					when "110010100111111" => rgb <= "101111";
					when "110010101000000" => rgb <= "101111";
					when "110010101000001" => rgb <= "101111";
					when "110010101000010" => rgb <= "101111";
					when "110010101000011" => rgb <= "101111";
					when "110010101000100" => rgb <= "101111";
					when "110010101000101" => rgb <= "101111";
					when "110010101000110" => rgb <= "101111";
					when "110010101000111" => rgb <= "101111";
					when "110010101001000" => rgb <= "101111";
					when "110010101001001" => rgb <= "101111";
					when "110010101001010" => rgb <= "101111";
					when "110010101001011" => rgb <= "101111";
					when "110010101001100" => rgb <= "101111";
					when "110010101001101" => rgb <= "101111";
					when "110010101001110" => rgb <= "101111";
					when "110010101001111" => rgb <= "101111";
					when "110010101010000" => rgb <= "101111";
					when "110010101010001" => rgb <= "101111";
					when "110010101010010" => rgb <= "101111";
					when "110010101010011" => rgb <= "101111";
					when "110010101010100" => rgb <= "101111";
					when "110010101010101" => rgb <= "101111";
					when "110010101010110" => rgb <= "101111";
					when "110010101010111" => rgb <= "101111";
					when "110010101011000" => rgb <= "101111";
					when "110010101011001" => rgb <= "101111";
					when "110010101011010" => rgb <= "101111";
					when "110010101011011" => rgb <= "101111";
					when "110010101011100" => rgb <= "101111";
					when "110010101011101" => rgb <= "101111";
					when "110010101011110" => rgb <= "101111";
					when "110010101011111" => rgb <= "101111";
					when "110010101100000" => rgb <= "101111";
					when "110010101100001" => rgb <= "101111";
					when "110010101100010" => rgb <= "101111";
					when "110010101100011" => rgb <= "101111";
					when "110010101100100" => rgb <= "101111";
					when "110010101100101" => rgb <= "101111";
					when "110010101100110" => rgb <= "101111";
					when "110010101100111" => rgb <= "101111";
					when "110010101101000" => rgb <= "101111";
					when "110010101101001" => rgb <= "101111";
					when "110010101101010" => rgb <= "101111";
					when "110010101101011" => rgb <= "101111";
					when "110010101101100" => rgb <= "101111";
					when "110010101101101" => rgb <= "101111";
					when "110010101101110" => rgb <= "101111";
					when "110010101101111" => rgb <= "101111";
					when "110010101110000" => rgb <= "101111";
					when "110010101110001" => rgb <= "101111";
					when "110010101110010" => rgb <= "101111";
					when "110010101110011" => rgb <= "101111";
					when "110010101110100" => rgb <= "101111";
					when "110010101110101" => rgb <= "101111";
					when "110010101110110" => rgb <= "101111";
					when "110010101110111" => rgb <= "101111";
					when "110010101111000" => rgb <= "101111";
					when "110010101111001" => rgb <= "101111";
					when "110010101111010" => rgb <= "101111";
					when "110010101111011" => rgb <= "101111";
					when "110010101111100" => rgb <= "101111";
					when "110010101111101" => rgb <= "101111";
					when "110010101111110" => rgb <= "101111";
					when "110010101111111" => rgb <= "101111";
					when "110010110000000" => rgb <= "101111";
					when "110010110000001" => rgb <= "101111";
					when "110010110000010" => rgb <= "101111";
					when "110010110000011" => rgb <= "101111";
					when "110010110000100" => rgb <= "101111";
					when "110010110000101" => rgb <= "101111";
					when "110010110000110" => rgb <= "101111";
					when "110010110000111" => rgb <= "101111";
					when "110010110001000" => rgb <= "101111";
					when "110010110001001" => rgb <= "101111";
					when "110010110001010" => rgb <= "000011";
					when "110010110001011" => rgb <= "000011";
					when "110010110001100" => rgb <= "101111";
					when "110010110001101" => rgb <= "101111";
					when "110010110001110" => rgb <= "101111";
					when "110010110001111" => rgb <= "101111";
					when "110010110010000" => rgb <= "101111";
					when "110010110010001" => rgb <= "101111";
					when "110010110010010" => rgb <= "101111";
					when "110010110010011" => rgb <= "101111";
					when "110010110010100" => rgb <= "101111";
					when "110010110010101" => rgb <= "101111";
					when "110010110010110" => rgb <= "101111";
					when "110010110010111" => rgb <= "101111";
					when "110010110011000" => rgb <= "101111";
					when "110010110011001" => rgb <= "101111";
					when "110010110011010" => rgb <= "101111";
					when "110010110011011" => rgb <= "101111";
					when "110010110011100" => rgb <= "101111";
					when "110010110011101" => rgb <= "101111";
					when "110010110011110" => rgb <= "101111";
					when "110010110011111" => rgb <= "101111";
					when "110011000000000" => rgb <= "101111";
					when "110011000000001" => rgb <= "101111";
					when "110011000000010" => rgb <= "101111";
					when "110011000000011" => rgb <= "101111";
					when "110011000000100" => rgb <= "101111";
					when "110011000000101" => rgb <= "101111";
					when "110011000000110" => rgb <= "101111";
					when "110011000000111" => rgb <= "101111";
					when "110011000001000" => rgb <= "101111";
					when "110011000001001" => rgb <= "101111";
					when "110011000001010" => rgb <= "101111";
					when "110011000001011" => rgb <= "101111";
					when "110011000001100" => rgb <= "101111";
					when "110011000001101" => rgb <= "101111";
					when "110011000001110" => rgb <= "101111";
					when "110011000001111" => rgb <= "101111";
					when "110011000010000" => rgb <= "101111";
					when "110011000010001" => rgb <= "101111";
					when "110011000010010" => rgb <= "101111";
					when "110011000010011" => rgb <= "101111";
					when "110011000010100" => rgb <= "101111";
					when "110011000010101" => rgb <= "101111";
					when "110011000010110" => rgb <= "101111";
					when "110011000010111" => rgb <= "101111";
					when "110011000011000" => rgb <= "101111";
					when "110011000011001" => rgb <= "101111";
					when "110011000011010" => rgb <= "101111";
					when "110011000011011" => rgb <= "101111";
					when "110011000011100" => rgb <= "101111";
					when "110011000011101" => rgb <= "101111";
					when "110011000011110" => rgb <= "000000";
					when "110011000011111" => rgb <= "000000";
					when "110011000100000" => rgb <= "100100";
					when "110011000100001" => rgb <= "100100";
					when "110011000100010" => rgb <= "100100";
					when "110011000100011" => rgb <= "100100";
					when "110011000100100" => rgb <= "100100";
					when "110011000100101" => rgb <= "100100";
					when "110011000100110" => rgb <= "100100";
					when "110011000100111" => rgb <= "100100";
					when "110011000101000" => rgb <= "100100";
					when "110011000101001" => rgb <= "100100";
					when "110011000101010" => rgb <= "100100";
					when "110011000101011" => rgb <= "100100";
					when "110011000101100" => rgb <= "100100";
					when "110011000101101" => rgb <= "100100";
					when "110011000101110" => rgb <= "100100";
					when "110011000101111" => rgb <= "100100";
					when "110011000110000" => rgb <= "100100";
					when "110011000110001" => rgb <= "100100";
					when "110011000110010" => rgb <= "100100";
					when "110011000110011" => rgb <= "100100";
					when "110011000110100" => rgb <= "010000";
					when "110011000110101" => rgb <= "010000";
					when "110011000110110" => rgb <= "000000";
					when "110011000110111" => rgb <= "000000";
					when "110011000111000" => rgb <= "000000";
					when "110011000111001" => rgb <= "000000";
					when "110011000111010" => rgb <= "101111";
					when "110011000111011" => rgb <= "101111";
					when "110011000111100" => rgb <= "101111";
					when "110011000111101" => rgb <= "101111";
					when "110011000111110" => rgb <= "101111";
					when "110011000111111" => rgb <= "101111";
					when "110011001000000" => rgb <= "101111";
					when "110011001000001" => rgb <= "101111";
					when "110011001000010" => rgb <= "101111";
					when "110011001000011" => rgb <= "101111";
					when "110011001000100" => rgb <= "101111";
					when "110011001000101" => rgb <= "101111";
					when "110011001000110" => rgb <= "101111";
					when "110011001000111" => rgb <= "101111";
					when "110011001001000" => rgb <= "101111";
					when "110011001001001" => rgb <= "101111";
					when "110011001001010" => rgb <= "101111";
					when "110011001001011" => rgb <= "101111";
					when "110011001001100" => rgb <= "101111";
					when "110011001001101" => rgb <= "101111";
					when "110011001001110" => rgb <= "101111";
					when "110011001001111" => rgb <= "101111";
					when "110011001010000" => rgb <= "101111";
					when "110011001010001" => rgb <= "101111";
					when "110011001010010" => rgb <= "101111";
					when "110011001010011" => rgb <= "101111";
					when "110011001010100" => rgb <= "101111";
					when "110011001010101" => rgb <= "101111";
					when "110011001010110" => rgb <= "101111";
					when "110011001010111" => rgb <= "101111";
					when "110011001011000" => rgb <= "101111";
					when "110011001011001" => rgb <= "101111";
					when "110011001011010" => rgb <= "101111";
					when "110011001011011" => rgb <= "101111";
					when "110011001011100" => rgb <= "101111";
					when "110011001011101" => rgb <= "101111";
					when "110011001011110" => rgb <= "101111";
					when "110011001011111" => rgb <= "101111";
					when "110011001100000" => rgb <= "101111";
					when "110011001100001" => rgb <= "101111";
					when "110011001100010" => rgb <= "101111";
					when "110011001100011" => rgb <= "101111";
					when "110011001100100" => rgb <= "101111";
					when "110011001100101" => rgb <= "101111";
					when "110011001100110" => rgb <= "101111";
					when "110011001100111" => rgb <= "101111";
					when "110011001101000" => rgb <= "101111";
					when "110011001101001" => rgb <= "101111";
					when "110011001101010" => rgb <= "101111";
					when "110011001101011" => rgb <= "101111";
					when "110011001101100" => rgb <= "101111";
					when "110011001101101" => rgb <= "101111";
					when "110011001101110" => rgb <= "101111";
					when "110011001101111" => rgb <= "101111";
					when "110011001110000" => rgb <= "101111";
					when "110011001110001" => rgb <= "101111";
					when "110011001110010" => rgb <= "101111";
					when "110011001110011" => rgb <= "101111";
					when "110011001110100" => rgb <= "101111";
					when "110011001110101" => rgb <= "101111";
					when "110011001110110" => rgb <= "101111";
					when "110011001110111" => rgb <= "101111";
					when "110011001111000" => rgb <= "101111";
					when "110011001111001" => rgb <= "101111";
					when "110011001111010" => rgb <= "101111";
					when "110011001111011" => rgb <= "101111";
					when "110011001111100" => rgb <= "101111";
					when "110011001111101" => rgb <= "101111";
					when "110011001111110" => rgb <= "101111";
					when "110011001111111" => rgb <= "101111";
					when "110011010000000" => rgb <= "101111";
					when "110011010000001" => rgb <= "101111";
					when "110011010000010" => rgb <= "101111";
					when "110011010000011" => rgb <= "101111";
					when "110011010000100" => rgb <= "101111";
					when "110011010000101" => rgb <= "101111";
					when "110011010000110" => rgb <= "101111";
					when "110011010000111" => rgb <= "101111";
					when "110011010001000" => rgb <= "101111";
					when "110011010001001" => rgb <= "101111";
					when "110011010001010" => rgb <= "101111";
					when "110011010001011" => rgb <= "101111";
					when "110011010001100" => rgb <= "101111";
					when "110011010001101" => rgb <= "101111";
					when "110011010001110" => rgb <= "101111";
					when "110011010001111" => rgb <= "101111";
					when "110011010010000" => rgb <= "101111";
					when "110011010010001" => rgb <= "101111";
					when "110011010010010" => rgb <= "101111";
					when "110011010010011" => rgb <= "101111";
					when "110011010010100" => rgb <= "101111";
					when "110011010010101" => rgb <= "101111";
					when "110011010010110" => rgb <= "101111";
					when "110011010010111" => rgb <= "101111";
					when "110011010011000" => rgb <= "101111";
					when "110011010011001" => rgb <= "101111";
					when "110011010011010" => rgb <= "101111";
					when "110011010011011" => rgb <= "101111";
					when "110011010011100" => rgb <= "101111";
					when "110011010011101" => rgb <= "101111";
					when "110011010011110" => rgb <= "101111";
					when "110011010011111" => rgb <= "101111";
					when "110011100000000" => rgb <= "101111";
					when "110011100000001" => rgb <= "101111";
					when "110011100000010" => rgb <= "101111";
					when "110011100000011" => rgb <= "101111";
					when "110011100000100" => rgb <= "101111";
					when "110011100000101" => rgb <= "101111";
					when "110011100000110" => rgb <= "101111";
					when "110011100000111" => rgb <= "101111";
					when "110011100001000" => rgb <= "101111";
					when "110011100001001" => rgb <= "101111";
					when "110011100001010" => rgb <= "101111";
					when "110011100001011" => rgb <= "101111";
					when "110011100001100" => rgb <= "101111";
					when "110011100001101" => rgb <= "101111";
					when "110011100001110" => rgb <= "101111";
					when "110011100001111" => rgb <= "101111";
					when "110011100010000" => rgb <= "101111";
					when "110011100010001" => rgb <= "101111";
					when "110011100010010" => rgb <= "101111";
					when "110011100010011" => rgb <= "101111";
					when "110011100010100" => rgb <= "101111";
					when "110011100010101" => rgb <= "101111";
					when "110011100010110" => rgb <= "101111";
					when "110011100010111" => rgb <= "101111";
					when "110011100011000" => rgb <= "101111";
					when "110011100011001" => rgb <= "101111";
					when "110011100011010" => rgb <= "101111";
					when "110011100011011" => rgb <= "101111";
					when "110011100011100" => rgb <= "101111";
					when "110011100011101" => rgb <= "101111";
					when "110011100011110" => rgb <= "000000";
					when "110011100011111" => rgb <= "000000";
					when "110011100100000" => rgb <= "100100";
					when "110011100100001" => rgb <= "100100";
					when "110011100100010" => rgb <= "100100";
					when "110011100100011" => rgb <= "100100";
					when "110011100100100" => rgb <= "100100";
					when "110011100100101" => rgb <= "100100";
					when "110011100100110" => rgb <= "100100";
					when "110011100100111" => rgb <= "100100";
					when "110011100101000" => rgb <= "100100";
					when "110011100101001" => rgb <= "100100";
					when "110011100101010" => rgb <= "100100";
					when "110011100101011" => rgb <= "100100";
					when "110011100101100" => rgb <= "100100";
					when "110011100101101" => rgb <= "100100";
					when "110011100101110" => rgb <= "100100";
					when "110011100101111" => rgb <= "100100";
					when "110011100110000" => rgb <= "100100";
					when "110011100110001" => rgb <= "100100";
					when "110011100110010" => rgb <= "100100";
					when "110011100110011" => rgb <= "100100";
					when "110011100110100" => rgb <= "010000";
					when "110011100110101" => rgb <= "010000";
					when "110011100110110" => rgb <= "000000";
					when "110011100110111" => rgb <= "000000";
					when "110011100111000" => rgb <= "000000";
					when "110011100111001" => rgb <= "000000";
					when "110011100111010" => rgb <= "101111";
					when "110011100111011" => rgb <= "101111";
					when "110011100111100" => rgb <= "101111";
					when "110011100111101" => rgb <= "101111";
					when "110011100111110" => rgb <= "101111";
					when "110011100111111" => rgb <= "101111";
					when "110011101000000" => rgb <= "101111";
					when "110011101000001" => rgb <= "101111";
					when "110011101000010" => rgb <= "101111";
					when "110011101000011" => rgb <= "101111";
					when "110011101000100" => rgb <= "101111";
					when "110011101000101" => rgb <= "101111";
					when "110011101000110" => rgb <= "101111";
					when "110011101000111" => rgb <= "101111";
					when "110011101001000" => rgb <= "101111";
					when "110011101001001" => rgb <= "101111";
					when "110011101001010" => rgb <= "101111";
					when "110011101001011" => rgb <= "101111";
					when "110011101001100" => rgb <= "101111";
					when "110011101001101" => rgb <= "101111";
					when "110011101001110" => rgb <= "101111";
					when "110011101001111" => rgb <= "101111";
					when "110011101010000" => rgb <= "101111";
					when "110011101010001" => rgb <= "101111";
					when "110011101010010" => rgb <= "101111";
					when "110011101010011" => rgb <= "101111";
					when "110011101010100" => rgb <= "101111";
					when "110011101010101" => rgb <= "101111";
					when "110011101010110" => rgb <= "101111";
					when "110011101010111" => rgb <= "101111";
					when "110011101011000" => rgb <= "101111";
					when "110011101011001" => rgb <= "101111";
					when "110011101011010" => rgb <= "101111";
					when "110011101011011" => rgb <= "101111";
					when "110011101011100" => rgb <= "101111";
					when "110011101011101" => rgb <= "101111";
					when "110011101011110" => rgb <= "101111";
					when "110011101011111" => rgb <= "101111";
					when "110011101100000" => rgb <= "101111";
					when "110011101100001" => rgb <= "101111";
					when "110011101100010" => rgb <= "101111";
					when "110011101100011" => rgb <= "101111";
					when "110011101100100" => rgb <= "101111";
					when "110011101100101" => rgb <= "101111";
					when "110011101100110" => rgb <= "101111";
					when "110011101100111" => rgb <= "101111";
					when "110011101101000" => rgb <= "101111";
					when "110011101101001" => rgb <= "101111";
					when "110011101101010" => rgb <= "101111";
					when "110011101101011" => rgb <= "101111";
					when "110011101101100" => rgb <= "101111";
					when "110011101101101" => rgb <= "101111";
					when "110011101101110" => rgb <= "101111";
					when "110011101101111" => rgb <= "101111";
					when "110011101110000" => rgb <= "101111";
					when "110011101110001" => rgb <= "101111";
					when "110011101110010" => rgb <= "101111";
					when "110011101110011" => rgb <= "101111";
					when "110011101110100" => rgb <= "101111";
					when "110011101110101" => rgb <= "101111";
					when "110011101110110" => rgb <= "101111";
					when "110011101110111" => rgb <= "101111";
					when "110011101111000" => rgb <= "101111";
					when "110011101111001" => rgb <= "101111";
					when "110011101111010" => rgb <= "101111";
					when "110011101111011" => rgb <= "101111";
					when "110011101111100" => rgb <= "101111";
					when "110011101111101" => rgb <= "101111";
					when "110011101111110" => rgb <= "101111";
					when "110011101111111" => rgb <= "101111";
					when "110011110000000" => rgb <= "101111";
					when "110011110000001" => rgb <= "101111";
					when "110011110000010" => rgb <= "101111";
					when "110011110000011" => rgb <= "101111";
					when "110011110000100" => rgb <= "101111";
					when "110011110000101" => rgb <= "101111";
					when "110011110000110" => rgb <= "101111";
					when "110011110000111" => rgb <= "101111";
					when "110011110001000" => rgb <= "101111";
					when "110011110001001" => rgb <= "101111";
					when "110011110001010" => rgb <= "101111";
					when "110011110001011" => rgb <= "101111";
					when "110011110001100" => rgb <= "101111";
					when "110011110001101" => rgb <= "101111";
					when "110011110001110" => rgb <= "101111";
					when "110011110001111" => rgb <= "101111";
					when "110011110010000" => rgb <= "101111";
					when "110011110010001" => rgb <= "101111";
					when "110011110010010" => rgb <= "101111";
					when "110011110010011" => rgb <= "101111";
					when "110011110010100" => rgb <= "101111";
					when "110011110010101" => rgb <= "101111";
					when "110011110010110" => rgb <= "101111";
					when "110011110010111" => rgb <= "101111";
					when "110011110011000" => rgb <= "101111";
					when "110011110011001" => rgb <= "101111";
					when "110011110011010" => rgb <= "101111";
					when "110011110011011" => rgb <= "101111";
					when "110011110011100" => rgb <= "101111";
					when "110011110011101" => rgb <= "101111";
					when "110011110011110" => rgb <= "101111";
					when "110011110011111" => rgb <= "101111";
					when "110100000000000" => rgb <= "101111";
					when "110100000000001" => rgb <= "101111";
					when "110100000000010" => rgb <= "101111";
					when "110100000000011" => rgb <= "101111";
					when "110100000000100" => rgb <= "101111";
					when "110100000000101" => rgb <= "101111";
					when "110100000000110" => rgb <= "101111";
					when "110100000000111" => rgb <= "101111";
					when "110100000001000" => rgb <= "101111";
					when "110100000001001" => rgb <= "101111";
					when "110100000001010" => rgb <= "101111";
					when "110100000001011" => rgb <= "101111";
					when "110100000001100" => rgb <= "101111";
					when "110100000001101" => rgb <= "101111";
					when "110100000001110" => rgb <= "101111";
					when "110100000001111" => rgb <= "101111";
					when "110100000010000" => rgb <= "101111";
					when "110100000010001" => rgb <= "101111";
					when "110100000010010" => rgb <= "101111";
					when "110100000010011" => rgb <= "101111";
					when "110100000010100" => rgb <= "101111";
					when "110100000010101" => rgb <= "101111";
					when "110100000010110" => rgb <= "101111";
					when "110100000010111" => rgb <= "101111";
					when "110100000011000" => rgb <= "101111";
					when "110100000011001" => rgb <= "101111";
					when "110100000011010" => rgb <= "101111";
					when "110100000011011" => rgb <= "101111";
					when "110100000011100" => rgb <= "101111";
					when "110100000011101" => rgb <= "101111";
					when "110100000011110" => rgb <= "000000";
					when "110100000011111" => rgb <= "000000";
					when "110100000100000" => rgb <= "100100";
					when "110100000100001" => rgb <= "100100";
					when "110100000100010" => rgb <= "100100";
					when "110100000100011" => rgb <= "100100";
					when "110100000100100" => rgb <= "100100";
					when "110100000100101" => rgb <= "100100";
					when "110100000100110" => rgb <= "100100";
					when "110100000100111" => rgb <= "100100";
					when "110100000101000" => rgb <= "100100";
					when "110100000101001" => rgb <= "100100";
					when "110100000101010" => rgb <= "100100";
					when "110100000101011" => rgb <= "100100";
					when "110100000101100" => rgb <= "100100";
					when "110100000101101" => rgb <= "100100";
					when "110100000101110" => rgb <= "100100";
					when "110100000101111" => rgb <= "100100";
					when "110100000110000" => rgb <= "100100";
					when "110100000110001" => rgb <= "100100";
					when "110100000110010" => rgb <= "100100";
					when "110100000110011" => rgb <= "100100";
					when "110100000110100" => rgb <= "100100";
					when "110100000110101" => rgb <= "100100";
					when "110100000110110" => rgb <= "010000";
					when "110100000110111" => rgb <= "010000";
					when "110100000111000" => rgb <= "000000";
					when "110100000111001" => rgb <= "000000";
					when "110100000111010" => rgb <= "101111";
					when "110100000111011" => rgb <= "101111";
					when "110100000111100" => rgb <= "101111";
					when "110100000111101" => rgb <= "101111";
					when "110100000111110" => rgb <= "101111";
					when "110100000111111" => rgb <= "101111";
					when "110100001000000" => rgb <= "101111";
					when "110100001000001" => rgb <= "101111";
					when "110100001000010" => rgb <= "101111";
					when "110100001000011" => rgb <= "101111";
					when "110100001000100" => rgb <= "101111";
					when "110100001000101" => rgb <= "101111";
					when "110100001000110" => rgb <= "101111";
					when "110100001000111" => rgb <= "101111";
					when "110100001001000" => rgb <= "101111";
					when "110100001001001" => rgb <= "101111";
					when "110100001001010" => rgb <= "101111";
					when "110100001001011" => rgb <= "101111";
					when "110100001001100" => rgb <= "101111";
					when "110100001001101" => rgb <= "101111";
					when "110100001001110" => rgb <= "101111";
					when "110100001001111" => rgb <= "101111";
					when "110100001010000" => rgb <= "101111";
					when "110100001010001" => rgb <= "101111";
					when "110100001010010" => rgb <= "101111";
					when "110100001010011" => rgb <= "101111";
					when "110100001010100" => rgb <= "101111";
					when "110100001010101" => rgb <= "101111";
					when "110100001010110" => rgb <= "101111";
					when "110100001010111" => rgb <= "101111";
					when "110100001011000" => rgb <= "101111";
					when "110100001011001" => rgb <= "101111";
					when "110100001011010" => rgb <= "101111";
					when "110100001011011" => rgb <= "101111";
					when "110100001011100" => rgb <= "101111";
					when "110100001011101" => rgb <= "101111";
					when "110100001011110" => rgb <= "101111";
					when "110100001011111" => rgb <= "101111";
					when "110100001100000" => rgb <= "101111";
					when "110100001100001" => rgb <= "101111";
					when "110100001100010" => rgb <= "101111";
					when "110100001100011" => rgb <= "101111";
					when "110100001100100" => rgb <= "101111";
					when "110100001100101" => rgb <= "101111";
					when "110100001100110" => rgb <= "101111";
					when "110100001100111" => rgb <= "101111";
					when "110100001101000" => rgb <= "101111";
					when "110100001101001" => rgb <= "101111";
					when "110100001101010" => rgb <= "101111";
					when "110100001101011" => rgb <= "101111";
					when "110100001101100" => rgb <= "101111";
					when "110100001101101" => rgb <= "101111";
					when "110100001101110" => rgb <= "101111";
					when "110100001101111" => rgb <= "101111";
					when "110100001110000" => rgb <= "101111";
					when "110100001110001" => rgb <= "101111";
					when "110100001110010" => rgb <= "101111";
					when "110100001110011" => rgb <= "101111";
					when "110100001110100" => rgb <= "101111";
					when "110100001110101" => rgb <= "101111";
					when "110100001110110" => rgb <= "101111";
					when "110100001110111" => rgb <= "101111";
					when "110100001111000" => rgb <= "101111";
					when "110100001111001" => rgb <= "101111";
					when "110100001111010" => rgb <= "101111";
					when "110100001111011" => rgb <= "101111";
					when "110100001111100" => rgb <= "101111";
					when "110100001111101" => rgb <= "101111";
					when "110100001111110" => rgb <= "101111";
					when "110100001111111" => rgb <= "101111";
					when "110100010000000" => rgb <= "101111";
					when "110100010000001" => rgb <= "101111";
					when "110100010000010" => rgb <= "101111";
					when "110100010000011" => rgb <= "101111";
					when "110100010000100" => rgb <= "101111";
					when "110100010000101" => rgb <= "101111";
					when "110100010000110" => rgb <= "101111";
					when "110100010000111" => rgb <= "101111";
					when "110100010001000" => rgb <= "101111";
					when "110100010001001" => rgb <= "101111";
					when "110100010001010" => rgb <= "101111";
					when "110100010001011" => rgb <= "101111";
					when "110100010001100" => rgb <= "101111";
					when "110100010001101" => rgb <= "101111";
					when "110100010001110" => rgb <= "101111";
					when "110100010001111" => rgb <= "101111";
					when "110100010010000" => rgb <= "101111";
					when "110100010010001" => rgb <= "101111";
					when "110100010010010" => rgb <= "101111";
					when "110100010010011" => rgb <= "101111";
					when "110100010010100" => rgb <= "101111";
					when "110100010010101" => rgb <= "101111";
					when "110100010010110" => rgb <= "101111";
					when "110100010010111" => rgb <= "101111";
					when "110100010011000" => rgb <= "101111";
					when "110100010011001" => rgb <= "101111";
					when "110100010011010" => rgb <= "101111";
					when "110100010011011" => rgb <= "101111";
					when "110100010011100" => rgb <= "101111";
					when "110100010011101" => rgb <= "101111";
					when "110100010011110" => rgb <= "101111";
					when "110100010011111" => rgb <= "101111";
					when "110100100000000" => rgb <= "101111";
					when "110100100000001" => rgb <= "101111";
					when "110100100000010" => rgb <= "101111";
					when "110100100000011" => rgb <= "101111";
					when "110100100000100" => rgb <= "101111";
					when "110100100000101" => rgb <= "101111";
					when "110100100000110" => rgb <= "101111";
					when "110100100000111" => rgb <= "101111";
					when "110100100001000" => rgb <= "101111";
					when "110100100001001" => rgb <= "101111";
					when "110100100001010" => rgb <= "101111";
					when "110100100001011" => rgb <= "101111";
					when "110100100001100" => rgb <= "101111";
					when "110100100001101" => rgb <= "101111";
					when "110100100001110" => rgb <= "101111";
					when "110100100001111" => rgb <= "101111";
					when "110100100010000" => rgb <= "101111";
					when "110100100010001" => rgb <= "101111";
					when "110100100010010" => rgb <= "101111";
					when "110100100010011" => rgb <= "101111";
					when "110100100010100" => rgb <= "101111";
					when "110100100010101" => rgb <= "101111";
					when "110100100010110" => rgb <= "101111";
					when "110100100010111" => rgb <= "101111";
					when "110100100011000" => rgb <= "101111";
					when "110100100011001" => rgb <= "101111";
					when "110100100011010" => rgb <= "101111";
					when "110100100011011" => rgb <= "101111";
					when "110100100011100" => rgb <= "101111";
					when "110100100011101" => rgb <= "101111";
					when "110100100011110" => rgb <= "000000";
					when "110100100011111" => rgb <= "000000";
					when "110100100100000" => rgb <= "100100";
					when "110100100100001" => rgb <= "100100";
					when "110100100100010" => rgb <= "100100";
					when "110100100100011" => rgb <= "100100";
					when "110100100100100" => rgb <= "100100";
					when "110100100100101" => rgb <= "100100";
					when "110100100100110" => rgb <= "100100";
					when "110100100100111" => rgb <= "100100";
					when "110100100101000" => rgb <= "100100";
					when "110100100101001" => rgb <= "100100";
					when "110100100101010" => rgb <= "100100";
					when "110100100101011" => rgb <= "100100";
					when "110100100101100" => rgb <= "100100";
					when "110100100101101" => rgb <= "100100";
					when "110100100101110" => rgb <= "100100";
					when "110100100101111" => rgb <= "100100";
					when "110100100110000" => rgb <= "100100";
					when "110100100110001" => rgb <= "100100";
					when "110100100110010" => rgb <= "100100";
					when "110100100110011" => rgb <= "100100";
					when "110100100110100" => rgb <= "100100";
					when "110100100110101" => rgb <= "100100";
					when "110100100110110" => rgb <= "010000";
					when "110100100110111" => rgb <= "010000";
					when "110100100111000" => rgb <= "000000";
					when "110100100111001" => rgb <= "000000";
					when "110100100111010" => rgb <= "101111";
					when "110100100111011" => rgb <= "101111";
					when "110100100111100" => rgb <= "101111";
					when "110100100111101" => rgb <= "101111";
					when "110100100111110" => rgb <= "101111";
					when "110100100111111" => rgb <= "101111";
					when "110100101000000" => rgb <= "101111";
					when "110100101000001" => rgb <= "101111";
					when "110100101000010" => rgb <= "101111";
					when "110100101000011" => rgb <= "101111";
					when "110100101000100" => rgb <= "101111";
					when "110100101000101" => rgb <= "101111";
					when "110100101000110" => rgb <= "101111";
					when "110100101000111" => rgb <= "101111";
					when "110100101001000" => rgb <= "101111";
					when "110100101001001" => rgb <= "101111";
					when "110100101001010" => rgb <= "101111";
					when "110100101001011" => rgb <= "101111";
					when "110100101001100" => rgb <= "101111";
					when "110100101001101" => rgb <= "101111";
					when "110100101001110" => rgb <= "101111";
					when "110100101001111" => rgb <= "101111";
					when "110100101010000" => rgb <= "101111";
					when "110100101010001" => rgb <= "101111";
					when "110100101010010" => rgb <= "101111";
					when "110100101010011" => rgb <= "101111";
					when "110100101010100" => rgb <= "101111";
					when "110100101010101" => rgb <= "101111";
					when "110100101010110" => rgb <= "101111";
					when "110100101010111" => rgb <= "101111";
					when "110100101011000" => rgb <= "101111";
					when "110100101011001" => rgb <= "101111";
					when "110100101011010" => rgb <= "101111";
					when "110100101011011" => rgb <= "101111";
					when "110100101011100" => rgb <= "101111";
					when "110100101011101" => rgb <= "101111";
					when "110100101011110" => rgb <= "101111";
					when "110100101011111" => rgb <= "101111";
					when "110100101100000" => rgb <= "101111";
					when "110100101100001" => rgb <= "101111";
					when "110100101100010" => rgb <= "101111";
					when "110100101100011" => rgb <= "101111";
					when "110100101100100" => rgb <= "101111";
					when "110100101100101" => rgb <= "101111";
					when "110100101100110" => rgb <= "101111";
					when "110100101100111" => rgb <= "101111";
					when "110100101101000" => rgb <= "101111";
					when "110100101101001" => rgb <= "101111";
					when "110100101101010" => rgb <= "101111";
					when "110100101101011" => rgb <= "101111";
					when "110100101101100" => rgb <= "101111";
					when "110100101101101" => rgb <= "101111";
					when "110100101101110" => rgb <= "101111";
					when "110100101101111" => rgb <= "101111";
					when "110100101110000" => rgb <= "101111";
					when "110100101110001" => rgb <= "101111";
					when "110100101110010" => rgb <= "101111";
					when "110100101110011" => rgb <= "101111";
					when "110100101110100" => rgb <= "101111";
					when "110100101110101" => rgb <= "101111";
					when "110100101110110" => rgb <= "101111";
					when "110100101110111" => rgb <= "101111";
					when "110100101111000" => rgb <= "101111";
					when "110100101111001" => rgb <= "101111";
					when "110100101111010" => rgb <= "101111";
					when "110100101111011" => rgb <= "101111";
					when "110100101111100" => rgb <= "101111";
					when "110100101111101" => rgb <= "101111";
					when "110100101111110" => rgb <= "101111";
					when "110100101111111" => rgb <= "101111";
					when "110100110000000" => rgb <= "101111";
					when "110100110000001" => rgb <= "101111";
					when "110100110000010" => rgb <= "101111";
					when "110100110000011" => rgb <= "101111";
					when "110100110000100" => rgb <= "101111";
					when "110100110000101" => rgb <= "101111";
					when "110100110000110" => rgb <= "101111";
					when "110100110000111" => rgb <= "101111";
					when "110100110001000" => rgb <= "101111";
					when "110100110001001" => rgb <= "101111";
					when "110100110001010" => rgb <= "101111";
					when "110100110001011" => rgb <= "101111";
					when "110100110001100" => rgb <= "101111";
					when "110100110001101" => rgb <= "101111";
					when "110100110001110" => rgb <= "101111";
					when "110100110001111" => rgb <= "101111";
					when "110100110010000" => rgb <= "101111";
					when "110100110010001" => rgb <= "101111";
					when "110100110010010" => rgb <= "101111";
					when "110100110010011" => rgb <= "101111";
					when "110100110010100" => rgb <= "101111";
					when "110100110010101" => rgb <= "101111";
					when "110100110010110" => rgb <= "101111";
					when "110100110010111" => rgb <= "101111";
					when "110100110011000" => rgb <= "101111";
					when "110100110011001" => rgb <= "101111";
					when "110100110011010" => rgb <= "101111";
					when "110100110011011" => rgb <= "101111";
					when "110100110011100" => rgb <= "101111";
					when "110100110011101" => rgb <= "101111";
					when "110100110011110" => rgb <= "101111";
					when "110100110011111" => rgb <= "101111";
					when "110101000000000" => rgb <= "101111";
					when "110101000000001" => rgb <= "101111";
					when "110101000000010" => rgb <= "101111";
					when "110101000000011" => rgb <= "101111";
					when "110101000000100" => rgb <= "101111";
					when "110101000000101" => rgb <= "101111";
					when "110101000000110" => rgb <= "101111";
					when "110101000000111" => rgb <= "101111";
					when "110101000001000" => rgb <= "101111";
					when "110101000001001" => rgb <= "101111";
					when "110101000001010" => rgb <= "101111";
					when "110101000001011" => rgb <= "101111";
					when "110101000001100" => rgb <= "101111";
					when "110101000001101" => rgb <= "101111";
					when "110101000001110" => rgb <= "101111";
					when "110101000001111" => rgb <= "101111";
					when "110101000010000" => rgb <= "101111";
					when "110101000010001" => rgb <= "101111";
					when "110101000010010" => rgb <= "101111";
					when "110101000010011" => rgb <= "101111";
					when "110101000010100" => rgb <= "101111";
					when "110101000010101" => rgb <= "101111";
					when "110101000010110" => rgb <= "101111";
					when "110101000010111" => rgb <= "101111";
					when "110101000011000" => rgb <= "101111";
					when "110101000011001" => rgb <= "101111";
					when "110101000011010" => rgb <= "101111";
					when "110101000011011" => rgb <= "101111";
					when "110101000011100" => rgb <= "000000";
					when "110101000011101" => rgb <= "000000";
					when "110101000011110" => rgb <= "100100";
					when "110101000011111" => rgb <= "100100";
					when "110101000100000" => rgb <= "100100";
					when "110101000100001" => rgb <= "100100";
					when "110101000100010" => rgb <= "100100";
					when "110101000100011" => rgb <= "100100";
					when "110101000100100" => rgb <= "100100";
					when "110101000100101" => rgb <= "100100";
					when "110101000100110" => rgb <= "100100";
					when "110101000100111" => rgb <= "100100";
					when "110101000101000" => rgb <= "100100";
					when "110101000101001" => rgb <= "100100";
					when "110101000101010" => rgb <= "100100";
					when "110101000101011" => rgb <= "100100";
					when "110101000101100" => rgb <= "100100";
					when "110101000101101" => rgb <= "100100";
					when "110101000101110" => rgb <= "100100";
					when "110101000101111" => rgb <= "100100";
					when "110101000110000" => rgb <= "100100";
					when "110101000110001" => rgb <= "100100";
					when "110101000110010" => rgb <= "100100";
					when "110101000110011" => rgb <= "100100";
					when "110101000110100" => rgb <= "100100";
					when "110101000110101" => rgb <= "100100";
					when "110101000110110" => rgb <= "100100";
					when "110101000110111" => rgb <= "100100";
					when "110101000111000" => rgb <= "010000";
					when "110101000111001" => rgb <= "010000";
					when "110101000111010" => rgb <= "000000";
					when "110101000111011" => rgb <= "000000";
					when "110101000111100" => rgb <= "101111";
					when "110101000111101" => rgb <= "101111";
					when "110101000111110" => rgb <= "101111";
					when "110101000111111" => rgb <= "101111";
					when "110101001000000" => rgb <= "101111";
					when "110101001000001" => rgb <= "101111";
					when "110101001000010" => rgb <= "101111";
					when "110101001000011" => rgb <= "101111";
					when "110101001000100" => rgb <= "101111";
					when "110101001000101" => rgb <= "101111";
					when "110101001000110" => rgb <= "101111";
					when "110101001000111" => rgb <= "101111";
					when "110101001001000" => rgb <= "101111";
					when "110101001001001" => rgb <= "101111";
					when "110101001001010" => rgb <= "101111";
					when "110101001001011" => rgb <= "101111";
					when "110101001001100" => rgb <= "101111";
					when "110101001001101" => rgb <= "101111";
					when "110101001001110" => rgb <= "101111";
					when "110101001001111" => rgb <= "101111";
					when "110101001010000" => rgb <= "101111";
					when "110101001010001" => rgb <= "101111";
					when "110101001010010" => rgb <= "101111";
					when "110101001010011" => rgb <= "101111";
					when "110101001010100" => rgb <= "101111";
					when "110101001010101" => rgb <= "101111";
					when "110101001010110" => rgb <= "101111";
					when "110101001010111" => rgb <= "101111";
					when "110101001011000" => rgb <= "101111";
					when "110101001011001" => rgb <= "101111";
					when "110101001011010" => rgb <= "101111";
					when "110101001011011" => rgb <= "101111";
					when "110101001011100" => rgb <= "101111";
					when "110101001011101" => rgb <= "101111";
					when "110101001011110" => rgb <= "101111";
					when "110101001011111" => rgb <= "101111";
					when "110101001100000" => rgb <= "101111";
					when "110101001100001" => rgb <= "101111";
					when "110101001100010" => rgb <= "101111";
					when "110101001100011" => rgb <= "101111";
					when "110101001100100" => rgb <= "101111";
					when "110101001100101" => rgb <= "101111";
					when "110101001100110" => rgb <= "101111";
					when "110101001100111" => rgb <= "101111";
					when "110101001101000" => rgb <= "101111";
					when "110101001101001" => rgb <= "101111";
					when "110101001101010" => rgb <= "101111";
					when "110101001101011" => rgb <= "101111";
					when "110101001101100" => rgb <= "101111";
					when "110101001101101" => rgb <= "101111";
					when "110101001101110" => rgb <= "101111";
					when "110101001101111" => rgb <= "101111";
					when "110101001110000" => rgb <= "101111";
					when "110101001110001" => rgb <= "101111";
					when "110101001110010" => rgb <= "101111";
					when "110101001110011" => rgb <= "101111";
					when "110101001110100" => rgb <= "101111";
					when "110101001110101" => rgb <= "101111";
					when "110101001110110" => rgb <= "101111";
					when "110101001110111" => rgb <= "101111";
					when "110101001111000" => rgb <= "101111";
					when "110101001111001" => rgb <= "101111";
					when "110101001111010" => rgb <= "101111";
					when "110101001111011" => rgb <= "101111";
					when "110101001111100" => rgb <= "101111";
					when "110101001111101" => rgb <= "101111";
					when "110101001111110" => rgb <= "101111";
					when "110101001111111" => rgb <= "101111";
					when "110101010000000" => rgb <= "101111";
					when "110101010000001" => rgb <= "101111";
					when "110101010000010" => rgb <= "101111";
					when "110101010000011" => rgb <= "101111";
					when "110101010000100" => rgb <= "101111";
					when "110101010000101" => rgb <= "101111";
					when "110101010000110" => rgb <= "101111";
					when "110101010000111" => rgb <= "101111";
					when "110101010001000" => rgb <= "101111";
					when "110101010001001" => rgb <= "101111";
					when "110101010001010" => rgb <= "101111";
					when "110101010001011" => rgb <= "101111";
					when "110101010001100" => rgb <= "101111";
					when "110101010001101" => rgb <= "101111";
					when "110101010001110" => rgb <= "101111";
					when "110101010001111" => rgb <= "101111";
					when "110101010010000" => rgb <= "101111";
					when "110101010010001" => rgb <= "101111";
					when "110101010010010" => rgb <= "101111";
					when "110101010010011" => rgb <= "101111";
					when "110101010010100" => rgb <= "101111";
					when "110101010010101" => rgb <= "101111";
					when "110101010010110" => rgb <= "101111";
					when "110101010010111" => rgb <= "101111";
					when "110101010011000" => rgb <= "101111";
					when "110101010011001" => rgb <= "101111";
					when "110101010011010" => rgb <= "101111";
					when "110101010011011" => rgb <= "101111";
					when "110101010011100" => rgb <= "101111";
					when "110101010011101" => rgb <= "101111";
					when "110101010011110" => rgb <= "101111";
					when "110101010011111" => rgb <= "101111";
					when "110101100000000" => rgb <= "101111";
					when "110101100000001" => rgb <= "101111";
					when "110101100000010" => rgb <= "101111";
					when "110101100000011" => rgb <= "101111";
					when "110101100000100" => rgb <= "101111";
					when "110101100000101" => rgb <= "101111";
					when "110101100000110" => rgb <= "101111";
					when "110101100000111" => rgb <= "101111";
					when "110101100001000" => rgb <= "101111";
					when "110101100001001" => rgb <= "101111";
					when "110101100001010" => rgb <= "101111";
					when "110101100001011" => rgb <= "101111";
					when "110101100001100" => rgb <= "101111";
					when "110101100001101" => rgb <= "101111";
					when "110101100001110" => rgb <= "101111";
					when "110101100001111" => rgb <= "101111";
					when "110101100010000" => rgb <= "101111";
					when "110101100010001" => rgb <= "101111";
					when "110101100010010" => rgb <= "101111";
					when "110101100010011" => rgb <= "101111";
					when "110101100010100" => rgb <= "101111";
					when "110101100010101" => rgb <= "101111";
					when "110101100010110" => rgb <= "101111";
					when "110101100010111" => rgb <= "101111";
					when "110101100011000" => rgb <= "101111";
					when "110101100011001" => rgb <= "101111";
					when "110101100011010" => rgb <= "101111";
					when "110101100011011" => rgb <= "101111";
					when "110101100011100" => rgb <= "000000";
					when "110101100011101" => rgb <= "000000";
					when "110101100011110" => rgb <= "100100";
					when "110101100011111" => rgb <= "100100";
					when "110101100100000" => rgb <= "100100";
					when "110101100100001" => rgb <= "100100";
					when "110101100100010" => rgb <= "100100";
					when "110101100100011" => rgb <= "100100";
					when "110101100100100" => rgb <= "100100";
					when "110101100100101" => rgb <= "100100";
					when "110101100100110" => rgb <= "100100";
					when "110101100100111" => rgb <= "100100";
					when "110101100101000" => rgb <= "100100";
					when "110101100101001" => rgb <= "100100";
					when "110101100101010" => rgb <= "100100";
					when "110101100101011" => rgb <= "100100";
					when "110101100101100" => rgb <= "100100";
					when "110101100101101" => rgb <= "100100";
					when "110101100101110" => rgb <= "100100";
					when "110101100101111" => rgb <= "100100";
					when "110101100110000" => rgb <= "100100";
					when "110101100110001" => rgb <= "100100";
					when "110101100110010" => rgb <= "100100";
					when "110101100110011" => rgb <= "100100";
					when "110101100110100" => rgb <= "100100";
					when "110101100110101" => rgb <= "100100";
					when "110101100110110" => rgb <= "100100";
					when "110101100110111" => rgb <= "100100";
					when "110101100111000" => rgb <= "010000";
					when "110101100111001" => rgb <= "010000";
					when "110101100111010" => rgb <= "000000";
					when "110101100111011" => rgb <= "000000";
					when "110101100111100" => rgb <= "101111";
					when "110101100111101" => rgb <= "101111";
					when "110101100111110" => rgb <= "101111";
					when "110101100111111" => rgb <= "101111";
					when "110101101000000" => rgb <= "101111";
					when "110101101000001" => rgb <= "101111";
					when "110101101000010" => rgb <= "101111";
					when "110101101000011" => rgb <= "101111";
					when "110101101000100" => rgb <= "101111";
					when "110101101000101" => rgb <= "101111";
					when "110101101000110" => rgb <= "101111";
					when "110101101000111" => rgb <= "101111";
					when "110101101001000" => rgb <= "101111";
					when "110101101001001" => rgb <= "101111";
					when "110101101001010" => rgb <= "101111";
					when "110101101001011" => rgb <= "101111";
					when "110101101001100" => rgb <= "101111";
					when "110101101001101" => rgb <= "101111";
					when "110101101001110" => rgb <= "101111";
					when "110101101001111" => rgb <= "101111";
					when "110101101010000" => rgb <= "101111";
					when "110101101010001" => rgb <= "101111";
					when "110101101010010" => rgb <= "101111";
					when "110101101010011" => rgb <= "101111";
					when "110101101010100" => rgb <= "101111";
					when "110101101010101" => rgb <= "101111";
					when "110101101010110" => rgb <= "101111";
					when "110101101010111" => rgb <= "101111";
					when "110101101011000" => rgb <= "101111";
					when "110101101011001" => rgb <= "101111";
					when "110101101011010" => rgb <= "101111";
					when "110101101011011" => rgb <= "101111";
					when "110101101011100" => rgb <= "101111";
					when "110101101011101" => rgb <= "101111";
					when "110101101011110" => rgb <= "101111";
					when "110101101011111" => rgb <= "101111";
					when "110101101100000" => rgb <= "101111";
					when "110101101100001" => rgb <= "101111";
					when "110101101100010" => rgb <= "101111";
					when "110101101100011" => rgb <= "101111";
					when "110101101100100" => rgb <= "101111";
					when "110101101100101" => rgb <= "101111";
					when "110101101100110" => rgb <= "101111";
					when "110101101100111" => rgb <= "101111";
					when "110101101101000" => rgb <= "101111";
					when "110101101101001" => rgb <= "101111";
					when "110101101101010" => rgb <= "101111";
					when "110101101101011" => rgb <= "101111";
					when "110101101101100" => rgb <= "101111";
					when "110101101101101" => rgb <= "101111";
					when "110101101101110" => rgb <= "101111";
					when "110101101101111" => rgb <= "101111";
					when "110101101110000" => rgb <= "101111";
					when "110101101110001" => rgb <= "101111";
					when "110101101110010" => rgb <= "101111";
					when "110101101110011" => rgb <= "101111";
					when "110101101110100" => rgb <= "101111";
					when "110101101110101" => rgb <= "101111";
					when "110101101110110" => rgb <= "101111";
					when "110101101110111" => rgb <= "101111";
					when "110101101111000" => rgb <= "101111";
					when "110101101111001" => rgb <= "101111";
					when "110101101111010" => rgb <= "101111";
					when "110101101111011" => rgb <= "101111";
					when "110101101111100" => rgb <= "101111";
					when "110101101111101" => rgb <= "101111";
					when "110101101111110" => rgb <= "101111";
					when "110101101111111" => rgb <= "101111";
					when "110101110000000" => rgb <= "101111";
					when "110101110000001" => rgb <= "101111";
					when "110101110000010" => rgb <= "101111";
					when "110101110000011" => rgb <= "101111";
					when "110101110000100" => rgb <= "101111";
					when "110101110000101" => rgb <= "101111";
					when "110101110000110" => rgb <= "101111";
					when "110101110000111" => rgb <= "101111";
					when "110101110001000" => rgb <= "101111";
					when "110101110001001" => rgb <= "101111";
					when "110101110001010" => rgb <= "101111";
					when "110101110001011" => rgb <= "101111";
					when "110101110001100" => rgb <= "101111";
					when "110101110001101" => rgb <= "101111";
					when "110101110001110" => rgb <= "101111";
					when "110101110001111" => rgb <= "101111";
					when "110101110010000" => rgb <= "101111";
					when "110101110010001" => rgb <= "101111";
					when "110101110010010" => rgb <= "101111";
					when "110101110010011" => rgb <= "101111";
					when "110101110010100" => rgb <= "101111";
					when "110101110010101" => rgb <= "101111";
					when "110101110010110" => rgb <= "101111";
					when "110101110010111" => rgb <= "101111";
					when "110101110011000" => rgb <= "101111";
					when "110101110011001" => rgb <= "101111";
					when "110101110011010" => rgb <= "101111";
					when "110101110011011" => rgb <= "101111";
					when "110101110011100" => rgb <= "101111";
					when "110101110011101" => rgb <= "101111";
					when "110101110011110" => rgb <= "101111";
					when "110101110011111" => rgb <= "101111";
					when "110110000000000" => rgb <= "101111";
					when "110110000000001" => rgb <= "101111";
					when "110110000000010" => rgb <= "101111";
					when "110110000000011" => rgb <= "101111";
					when "110110000000100" => rgb <= "101111";
					when "110110000000101" => rgb <= "101111";
					when "110110000000110" => rgb <= "101111";
					when "110110000000111" => rgb <= "101111";
					when "110110000001000" => rgb <= "101111";
					when "110110000001001" => rgb <= "101111";
					when "110110000001010" => rgb <= "101111";
					when "110110000001011" => rgb <= "101111";
					when "110110000001100" => rgb <= "101111";
					when "110110000001101" => rgb <= "101111";
					when "110110000001110" => rgb <= "101111";
					when "110110000001111" => rgb <= "101111";
					when "110110000010000" => rgb <= "101111";
					when "110110000010001" => rgb <= "101111";
					when "110110000010010" => rgb <= "101111";
					when "110110000010011" => rgb <= "101111";
					when "110110000010100" => rgb <= "101111";
					when "110110000010101" => rgb <= "101111";
					when "110110000010110" => rgb <= "101111";
					when "110110000010111" => rgb <= "101111";
					when "110110000011000" => rgb <= "101111";
					when "110110000011001" => rgb <= "101111";
					when "110110000011010" => rgb <= "101111";
					when "110110000011011" => rgb <= "101111";
					when "110110000011100" => rgb <= "000000";
					when "110110000011101" => rgb <= "000000";
					when "110110000011110" => rgb <= "100100";
					when "110110000011111" => rgb <= "100100";
					when "110110000100000" => rgb <= "100100";
					when "110110000100001" => rgb <= "100100";
					when "110110000100010" => rgb <= "100100";
					when "110110000100011" => rgb <= "100100";
					when "110110000100100" => rgb <= "100100";
					when "110110000100101" => rgb <= "100100";
					when "110110000100110" => rgb <= "100100";
					when "110110000100111" => rgb <= "100100";
					when "110110000101000" => rgb <= "100100";
					when "110110000101001" => rgb <= "100100";
					when "110110000101010" => rgb <= "100100";
					when "110110000101011" => rgb <= "100100";
					when "110110000101100" => rgb <= "100100";
					when "110110000101101" => rgb <= "100100";
					when "110110000101110" => rgb <= "100100";
					when "110110000101111" => rgb <= "100100";
					when "110110000110000" => rgb <= "100100";
					when "110110000110001" => rgb <= "100100";
					when "110110000110010" => rgb <= "100100";
					when "110110000110011" => rgb <= "100100";
					when "110110000110100" => rgb <= "100100";
					when "110110000110101" => rgb <= "100100";
					when "110110000110110" => rgb <= "100100";
					when "110110000110111" => rgb <= "100100";
					when "110110000111000" => rgb <= "010000";
					when "110110000111001" => rgb <= "010000";
					when "110110000111010" => rgb <= "000000";
					when "110110000111011" => rgb <= "000000";
					when "110110000111100" => rgb <= "101111";
					when "110110000111101" => rgb <= "101111";
					when "110110000111110" => rgb <= "101111";
					when "110110000111111" => rgb <= "101111";
					when "110110001000000" => rgb <= "101111";
					when "110110001000001" => rgb <= "101111";
					when "110110001000010" => rgb <= "101111";
					when "110110001000011" => rgb <= "101111";
					when "110110001000100" => rgb <= "101111";
					when "110110001000101" => rgb <= "101111";
					when "110110001000110" => rgb <= "101111";
					when "110110001000111" => rgb <= "101111";
					when "110110001001000" => rgb <= "101111";
					when "110110001001001" => rgb <= "101111";
					when "110110001001010" => rgb <= "101111";
					when "110110001001011" => rgb <= "101111";
					when "110110001001100" => rgb <= "101111";
					when "110110001001101" => rgb <= "101111";
					when "110110001001110" => rgb <= "101111";
					when "110110001001111" => rgb <= "101111";
					when "110110001010000" => rgb <= "101111";
					when "110110001010001" => rgb <= "101111";
					when "110110001010010" => rgb <= "101111";
					when "110110001010011" => rgb <= "101111";
					when "110110001010100" => rgb <= "101111";
					when "110110001010101" => rgb <= "101111";
					when "110110001010110" => rgb <= "101111";
					when "110110001010111" => rgb <= "101111";
					when "110110001011000" => rgb <= "101111";
					when "110110001011001" => rgb <= "101111";
					when "110110001011010" => rgb <= "101111";
					when "110110001011011" => rgb <= "101111";
					when "110110001011100" => rgb <= "101111";
					when "110110001011101" => rgb <= "101111";
					when "110110001011110" => rgb <= "101111";
					when "110110001011111" => rgb <= "101111";
					when "110110001100000" => rgb <= "101111";
					when "110110001100001" => rgb <= "101111";
					when "110110001100010" => rgb <= "101111";
					when "110110001100011" => rgb <= "101111";
					when "110110001100100" => rgb <= "101111";
					when "110110001100101" => rgb <= "101111";
					when "110110001100110" => rgb <= "101111";
					when "110110001100111" => rgb <= "101111";
					when "110110001101000" => rgb <= "101111";
					when "110110001101001" => rgb <= "101111";
					when "110110001101010" => rgb <= "101111";
					when "110110001101011" => rgb <= "101111";
					when "110110001101100" => rgb <= "101111";
					when "110110001101101" => rgb <= "101111";
					when "110110001101110" => rgb <= "101111";
					when "110110001101111" => rgb <= "101111";
					when "110110001110000" => rgb <= "101111";
					when "110110001110001" => rgb <= "101111";
					when "110110001110010" => rgb <= "101111";
					when "110110001110011" => rgb <= "101111";
					when "110110001110100" => rgb <= "101111";
					when "110110001110101" => rgb <= "101111";
					when "110110001110110" => rgb <= "101111";
					when "110110001110111" => rgb <= "101111";
					when "110110001111000" => rgb <= "101111";
					when "110110001111001" => rgb <= "101111";
					when "110110001111010" => rgb <= "101111";
					when "110110001111011" => rgb <= "101111";
					when "110110001111100" => rgb <= "101111";
					when "110110001111101" => rgb <= "101111";
					when "110110001111110" => rgb <= "101111";
					when "110110001111111" => rgb <= "101111";
					when "110110010000000" => rgb <= "101111";
					when "110110010000001" => rgb <= "101111";
					when "110110010000010" => rgb <= "101111";
					when "110110010000011" => rgb <= "101111";
					when "110110010000100" => rgb <= "101111";
					when "110110010000101" => rgb <= "101111";
					when "110110010000110" => rgb <= "101111";
					when "110110010000111" => rgb <= "101111";
					when "110110010001000" => rgb <= "101111";
					when "110110010001001" => rgb <= "101111";
					when "110110010001010" => rgb <= "101111";
					when "110110010001011" => rgb <= "101111";
					when "110110010001100" => rgb <= "101111";
					when "110110010001101" => rgb <= "101111";
					when "110110010001110" => rgb <= "101111";
					when "110110010001111" => rgb <= "101111";
					when "110110010010000" => rgb <= "101111";
					when "110110010010001" => rgb <= "101111";
					when "110110010010010" => rgb <= "101111";
					when "110110010010011" => rgb <= "101111";
					when "110110010010100" => rgb <= "101111";
					when "110110010010101" => rgb <= "101111";
					when "110110010010110" => rgb <= "101111";
					when "110110010010111" => rgb <= "101111";
					when "110110010011000" => rgb <= "101111";
					when "110110010011001" => rgb <= "101111";
					when "110110010011010" => rgb <= "101111";
					when "110110010011011" => rgb <= "101111";
					when "110110010011100" => rgb <= "101111";
					when "110110010011101" => rgb <= "101111";
					when "110110010011110" => rgb <= "101111";
					when "110110010011111" => rgb <= "101111";
					when "110110100000000" => rgb <= "101111";
					when "110110100000001" => rgb <= "101111";
					when "110110100000010" => rgb <= "101111";
					when "110110100000011" => rgb <= "101111";
					when "110110100000100" => rgb <= "101111";
					when "110110100000101" => rgb <= "101111";
					when "110110100000110" => rgb <= "101111";
					when "110110100000111" => rgb <= "101111";
					when "110110100001000" => rgb <= "101111";
					when "110110100001001" => rgb <= "101111";
					when "110110100001010" => rgb <= "101111";
					when "110110100001011" => rgb <= "101111";
					when "110110100001100" => rgb <= "101111";
					when "110110100001101" => rgb <= "101111";
					when "110110100001110" => rgb <= "101111";
					when "110110100001111" => rgb <= "101111";
					when "110110100010000" => rgb <= "101111";
					when "110110100010001" => rgb <= "101111";
					when "110110100010010" => rgb <= "101111";
					when "110110100010011" => rgb <= "101111";
					when "110110100010100" => rgb <= "101111";
					when "110110100010101" => rgb <= "101111";
					when "110110100010110" => rgb <= "101111";
					when "110110100010111" => rgb <= "101111";
					when "110110100011000" => rgb <= "101111";
					when "110110100011001" => rgb <= "101111";
					when "110110100011010" => rgb <= "101111";
					when "110110100011011" => rgb <= "101111";
					when "110110100011100" => rgb <= "000000";
					when "110110100011101" => rgb <= "000000";
					when "110110100011110" => rgb <= "100100";
					when "110110100011111" => rgb <= "100100";
					when "110110100100000" => rgb <= "100100";
					when "110110100100001" => rgb <= "100100";
					when "110110100100010" => rgb <= "100100";
					when "110110100100011" => rgb <= "100100";
					when "110110100100100" => rgb <= "100100";
					when "110110100100101" => rgb <= "100100";
					when "110110100100110" => rgb <= "100100";
					when "110110100100111" => rgb <= "100100";
					when "110110100101000" => rgb <= "100100";
					when "110110100101001" => rgb <= "100100";
					when "110110100101010" => rgb <= "100100";
					when "110110100101011" => rgb <= "100100";
					when "110110100101100" => rgb <= "100100";
					when "110110100101101" => rgb <= "100100";
					when "110110100101110" => rgb <= "100100";
					when "110110100101111" => rgb <= "100100";
					when "110110100110000" => rgb <= "100100";
					when "110110100110001" => rgb <= "100100";
					when "110110100110010" => rgb <= "100100";
					when "110110100110011" => rgb <= "100100";
					when "110110100110100" => rgb <= "100100";
					when "110110100110101" => rgb <= "100100";
					when "110110100110110" => rgb <= "100100";
					when "110110100110111" => rgb <= "100100";
					when "110110100111000" => rgb <= "010000";
					when "110110100111001" => rgb <= "010000";
					when "110110100111010" => rgb <= "000000";
					when "110110100111011" => rgb <= "000000";
					when "110110100111100" => rgb <= "101111";
					when "110110100111101" => rgb <= "101111";
					when "110110100111110" => rgb <= "101111";
					when "110110100111111" => rgb <= "101111";
					when "110110101000000" => rgb <= "101111";
					when "110110101000001" => rgb <= "101111";
					when "110110101000010" => rgb <= "101111";
					when "110110101000011" => rgb <= "101111";
					when "110110101000100" => rgb <= "101111";
					when "110110101000101" => rgb <= "101111";
					when "110110101000110" => rgb <= "101111";
					when "110110101000111" => rgb <= "101111";
					when "110110101001000" => rgb <= "101111";
					when "110110101001001" => rgb <= "101111";
					when "110110101001010" => rgb <= "101111";
					when "110110101001011" => rgb <= "101111";
					when "110110101001100" => rgb <= "101111";
					when "110110101001101" => rgb <= "101111";
					when "110110101001110" => rgb <= "101111";
					when "110110101001111" => rgb <= "101111";
					when "110110101010000" => rgb <= "101111";
					when "110110101010001" => rgb <= "101111";
					when "110110101010010" => rgb <= "101111";
					when "110110101010011" => rgb <= "101111";
					when "110110101010100" => rgb <= "101111";
					when "110110101010101" => rgb <= "101111";
					when "110110101010110" => rgb <= "101111";
					when "110110101010111" => rgb <= "101111";
					when "110110101011000" => rgb <= "101111";
					when "110110101011001" => rgb <= "101111";
					when "110110101011010" => rgb <= "101111";
					when "110110101011011" => rgb <= "101111";
					when "110110101011100" => rgb <= "101111";
					when "110110101011101" => rgb <= "101111";
					when "110110101011110" => rgb <= "101111";
					when "110110101011111" => rgb <= "101111";
					when "110110101100000" => rgb <= "101111";
					when "110110101100001" => rgb <= "101111";
					when "110110101100010" => rgb <= "101111";
					when "110110101100011" => rgb <= "101111";
					when "110110101100100" => rgb <= "101111";
					when "110110101100101" => rgb <= "101111";
					when "110110101100110" => rgb <= "101111";
					when "110110101100111" => rgb <= "101111";
					when "110110101101000" => rgb <= "101111";
					when "110110101101001" => rgb <= "101111";
					when "110110101101010" => rgb <= "101111";
					when "110110101101011" => rgb <= "101111";
					when "110110101101100" => rgb <= "101111";
					when "110110101101101" => rgb <= "101111";
					when "110110101101110" => rgb <= "101111";
					when "110110101101111" => rgb <= "101111";
					when "110110101110000" => rgb <= "101111";
					when "110110101110001" => rgb <= "101111";
					when "110110101110010" => rgb <= "101111";
					when "110110101110011" => rgb <= "101111";
					when "110110101110100" => rgb <= "101111";
					when "110110101110101" => rgb <= "101111";
					when "110110101110110" => rgb <= "101111";
					when "110110101110111" => rgb <= "101111";
					when "110110101111000" => rgb <= "101111";
					when "110110101111001" => rgb <= "101111";
					when "110110101111010" => rgb <= "101111";
					when "110110101111011" => rgb <= "101111";
					when "110110101111100" => rgb <= "101111";
					when "110110101111101" => rgb <= "101111";
					when "110110101111110" => rgb <= "101111";
					when "110110101111111" => rgb <= "101111";
					when "110110110000000" => rgb <= "101111";
					when "110110110000001" => rgb <= "101111";
					when "110110110000010" => rgb <= "101111";
					when "110110110000011" => rgb <= "101111";
					when "110110110000100" => rgb <= "101111";
					when "110110110000101" => rgb <= "101111";
					when "110110110000110" => rgb <= "101111";
					when "110110110000111" => rgb <= "101111";
					when "110110110001000" => rgb <= "101111";
					when "110110110001001" => rgb <= "101111";
					when "110110110001010" => rgb <= "101111";
					when "110110110001011" => rgb <= "101111";
					when "110110110001100" => rgb <= "101111";
					when "110110110001101" => rgb <= "101111";
					when "110110110001110" => rgb <= "101111";
					when "110110110001111" => rgb <= "101111";
					when "110110110010000" => rgb <= "101111";
					when "110110110010001" => rgb <= "101111";
					when "110110110010010" => rgb <= "101111";
					when "110110110010011" => rgb <= "101111";
					when "110110110010100" => rgb <= "101111";
					when "110110110010101" => rgb <= "101111";
					when "110110110010110" => rgb <= "101111";
					when "110110110010111" => rgb <= "101111";
					when "110110110011000" => rgb <= "101111";
					when "110110110011001" => rgb <= "101111";
					when "110110110011010" => rgb <= "101111";
					when "110110110011011" => rgb <= "101111";
					when "110110110011100" => rgb <= "101111";
					when "110110110011101" => rgb <= "101111";
					when "110110110011110" => rgb <= "101111";
					when "110110110011111" => rgb <= "101111";
					when "110111000000000" => rgb <= "101111";
					when "110111000000001" => rgb <= "101111";
					when "110111000000010" => rgb <= "101111";
					when "110111000000011" => rgb <= "101111";
					when "110111000000100" => rgb <= "101111";
					when "110111000000101" => rgb <= "101111";
					when "110111000000110" => rgb <= "101111";
					when "110111000000111" => rgb <= "101111";
					when "110111000001000" => rgb <= "101111";
					when "110111000001001" => rgb <= "101111";
					when "110111000001010" => rgb <= "101111";
					when "110111000001011" => rgb <= "101111";
					when "110111000001100" => rgb <= "101111";
					when "110111000001101" => rgb <= "101111";
					when "110111000001110" => rgb <= "101111";
					when "110111000001111" => rgb <= "101111";
					when "110111000010000" => rgb <= "101111";
					when "110111000010001" => rgb <= "101111";
					when "110111000010010" => rgb <= "101111";
					when "110111000010011" => rgb <= "101111";
					when "110111000010100" => rgb <= "101111";
					when "110111000010101" => rgb <= "101111";
					when "110111000010110" => rgb <= "101111";
					when "110111000010111" => rgb <= "101111";
					when "110111000011000" => rgb <= "101111";
					when "110111000011001" => rgb <= "101111";
					when "110111000011010" => rgb <= "000000";
					when "110111000011011" => rgb <= "000000";
					when "110111000011100" => rgb <= "000000";
					when "110111000011101" => rgb <= "000000";
					when "110111000011110" => rgb <= "100100";
					when "110111000011111" => rgb <= "100100";
					when "110111000100000" => rgb <= "100100";
					when "110111000100001" => rgb <= "100100";
					when "110111000100010" => rgb <= "100100";
					when "110111000100011" => rgb <= "100100";
					when "110111000100100" => rgb <= "100100";
					when "110111000100101" => rgb <= "100100";
					when "110111000100110" => rgb <= "100100";
					when "110111000100111" => rgb <= "100100";
					when "110111000101000" => rgb <= "100100";
					when "110111000101001" => rgb <= "100100";
					when "110111000101010" => rgb <= "100100";
					when "110111000101011" => rgb <= "100100";
					when "110111000101100" => rgb <= "100100";
					when "110111000101101" => rgb <= "100100";
					when "110111000101110" => rgb <= "100100";
					when "110111000101111" => rgb <= "100100";
					when "110111000110000" => rgb <= "100100";
					when "110111000110001" => rgb <= "100100";
					when "110111000110010" => rgb <= "100100";
					when "110111000110011" => rgb <= "100100";
					when "110111000110100" => rgb <= "100100";
					when "110111000110101" => rgb <= "100100";
					when "110111000110110" => rgb <= "100100";
					when "110111000110111" => rgb <= "100100";
					when "110111000111000" => rgb <= "010000";
					when "110111000111001" => rgb <= "010000";
					when "110111000111010" => rgb <= "000000";
					when "110111000111011" => rgb <= "000000";
					when "110111000111100" => rgb <= "101111";
					when "110111000111101" => rgb <= "101111";
					when "110111000111110" => rgb <= "101111";
					when "110111000111111" => rgb <= "101111";
					when "110111001000000" => rgb <= "101111";
					when "110111001000001" => rgb <= "101111";
					when "110111001000010" => rgb <= "101111";
					when "110111001000011" => rgb <= "101111";
					when "110111001000100" => rgb <= "101111";
					when "110111001000101" => rgb <= "101111";
					when "110111001000110" => rgb <= "101111";
					when "110111001000111" => rgb <= "101111";
					when "110111001001000" => rgb <= "101111";
					when "110111001001001" => rgb <= "101111";
					when "110111001001010" => rgb <= "101111";
					when "110111001001011" => rgb <= "101111";
					when "110111001001100" => rgb <= "101111";
					when "110111001001101" => rgb <= "101111";
					when "110111001001110" => rgb <= "101111";
					when "110111001001111" => rgb <= "101111";
					when "110111001010000" => rgb <= "101111";
					when "110111001010001" => rgb <= "101111";
					when "110111001010010" => rgb <= "101111";
					when "110111001010011" => rgb <= "101111";
					when "110111001010100" => rgb <= "101111";
					when "110111001010101" => rgb <= "101111";
					when "110111001010110" => rgb <= "101111";
					when "110111001010111" => rgb <= "101111";
					when "110111001011000" => rgb <= "101111";
					when "110111001011001" => rgb <= "101111";
					when "110111001011010" => rgb <= "101111";
					when "110111001011011" => rgb <= "101111";
					when "110111001011100" => rgb <= "101111";
					when "110111001011101" => rgb <= "101111";
					when "110111001011110" => rgb <= "101111";
					when "110111001011111" => rgb <= "101111";
					when "110111001100000" => rgb <= "101111";
					when "110111001100001" => rgb <= "101111";
					when "110111001100010" => rgb <= "101111";
					when "110111001100011" => rgb <= "101111";
					when "110111001100100" => rgb <= "101111";
					when "110111001100101" => rgb <= "101111";
					when "110111001100110" => rgb <= "101111";
					when "110111001100111" => rgb <= "101111";
					when "110111001101000" => rgb <= "101111";
					when "110111001101001" => rgb <= "101111";
					when "110111001101010" => rgb <= "101111";
					when "110111001101011" => rgb <= "101111";
					when "110111001101100" => rgb <= "101111";
					when "110111001101101" => rgb <= "101111";
					when "110111001101110" => rgb <= "101111";
					when "110111001101111" => rgb <= "101111";
					when "110111001110000" => rgb <= "101111";
					when "110111001110001" => rgb <= "101111";
					when "110111001110010" => rgb <= "101111";
					when "110111001110011" => rgb <= "101111";
					when "110111001110100" => rgb <= "101111";
					when "110111001110101" => rgb <= "101111";
					when "110111001110110" => rgb <= "101111";
					when "110111001110111" => rgb <= "101111";
					when "110111001111000" => rgb <= "101111";
					when "110111001111001" => rgb <= "101111";
					when "110111001111010" => rgb <= "101111";
					when "110111001111011" => rgb <= "101111";
					when "110111001111100" => rgb <= "101111";
					when "110111001111101" => rgb <= "101111";
					when "110111001111110" => rgb <= "101111";
					when "110111001111111" => rgb <= "101111";
					when "110111010000000" => rgb <= "101111";
					when "110111010000001" => rgb <= "101111";
					when "110111010000010" => rgb <= "101111";
					when "110111010000011" => rgb <= "101111";
					when "110111010000100" => rgb <= "101111";
					when "110111010000101" => rgb <= "101111";
					when "110111010000110" => rgb <= "101111";
					when "110111010000111" => rgb <= "101111";
					when "110111010001000" => rgb <= "101111";
					when "110111010001001" => rgb <= "101111";
					when "110111010001010" => rgb <= "101111";
					when "110111010001011" => rgb <= "101111";
					when "110111010001100" => rgb <= "101111";
					when "110111010001101" => rgb <= "101111";
					when "110111010001110" => rgb <= "101111";
					when "110111010001111" => rgb <= "101111";
					when "110111010010000" => rgb <= "101111";
					when "110111010010001" => rgb <= "101111";
					when "110111010010010" => rgb <= "101111";
					when "110111010010011" => rgb <= "101111";
					when "110111010010100" => rgb <= "101111";
					when "110111010010101" => rgb <= "101111";
					when "110111010010110" => rgb <= "101111";
					when "110111010010111" => rgb <= "101111";
					when "110111010011000" => rgb <= "101111";
					when "110111010011001" => rgb <= "101111";
					when "110111010011010" => rgb <= "101111";
					when "110111010011011" => rgb <= "101111";
					when "110111010011100" => rgb <= "101111";
					when "110111010011101" => rgb <= "101111";
					when "110111010011110" => rgb <= "101111";
					when "110111010011111" => rgb <= "101111";
					when "110111100000000" => rgb <= "101111";
					when "110111100000001" => rgb <= "101111";
					when "110111100000010" => rgb <= "101111";
					when "110111100000011" => rgb <= "101111";
					when "110111100000100" => rgb <= "101111";
					when "110111100000101" => rgb <= "101111";
					when "110111100000110" => rgb <= "101111";
					when "110111100000111" => rgb <= "101111";
					when "110111100001000" => rgb <= "101111";
					when "110111100001001" => rgb <= "101111";
					when "110111100001010" => rgb <= "101111";
					when "110111100001011" => rgb <= "101111";
					when "110111100001100" => rgb <= "101111";
					when "110111100001101" => rgb <= "101111";
					when "110111100001110" => rgb <= "101111";
					when "110111100001111" => rgb <= "101111";
					when "110111100010000" => rgb <= "101111";
					when "110111100010001" => rgb <= "101111";
					when "110111100010010" => rgb <= "101111";
					when "110111100010011" => rgb <= "101111";
					when "110111100010100" => rgb <= "101111";
					when "110111100010101" => rgb <= "101111";
					when "110111100010110" => rgb <= "101111";
					when "110111100010111" => rgb <= "101111";
					when "110111100011000" => rgb <= "101111";
					when "110111100011001" => rgb <= "101111";
					when "110111100011010" => rgb <= "000000";
					when "110111100011011" => rgb <= "000000";
					when "110111100011100" => rgb <= "000000";
					when "110111100011101" => rgb <= "000000";
					when "110111100011110" => rgb <= "100100";
					when "110111100011111" => rgb <= "100100";
					when "110111100100000" => rgb <= "100100";
					when "110111100100001" => rgb <= "100100";
					when "110111100100010" => rgb <= "100100";
					when "110111100100011" => rgb <= "100100";
					when "110111100100100" => rgb <= "100100";
					when "110111100100101" => rgb <= "100100";
					when "110111100100110" => rgb <= "100100";
					when "110111100100111" => rgb <= "100100";
					when "110111100101000" => rgb <= "100100";
					when "110111100101001" => rgb <= "100100";
					when "110111100101010" => rgb <= "100100";
					when "110111100101011" => rgb <= "100100";
					when "110111100101100" => rgb <= "100100";
					when "110111100101101" => rgb <= "100100";
					when "110111100101110" => rgb <= "100100";
					when "110111100101111" => rgb <= "100100";
					when "110111100110000" => rgb <= "100100";
					when "110111100110001" => rgb <= "100100";
					when "110111100110010" => rgb <= "100100";
					when "110111100110011" => rgb <= "100100";
					when "110111100110100" => rgb <= "100100";
					when "110111100110101" => rgb <= "100100";
					when "110111100110110" => rgb <= "100100";
					when "110111100110111" => rgb <= "100100";
					when "110111100111000" => rgb <= "010000";
					when "110111100111001" => rgb <= "010000";
					when "110111100111010" => rgb <= "000000";
					when "110111100111011" => rgb <= "000000";
					when "110111100111100" => rgb <= "101111";
					when "110111100111101" => rgb <= "101111";
					when "110111100111110" => rgb <= "101111";
					when "110111100111111" => rgb <= "101111";
					when "110111101000000" => rgb <= "101111";
					when "110111101000001" => rgb <= "101111";
					when "110111101000010" => rgb <= "101111";
					when "110111101000011" => rgb <= "101111";
					when "110111101000100" => rgb <= "101111";
					when "110111101000101" => rgb <= "101111";
					when "110111101000110" => rgb <= "101111";
					when "110111101000111" => rgb <= "101111";
					when "110111101001000" => rgb <= "101111";
					when "110111101001001" => rgb <= "101111";
					when "110111101001010" => rgb <= "101111";
					when "110111101001011" => rgb <= "101111";
					when "110111101001100" => rgb <= "101111";
					when "110111101001101" => rgb <= "101111";
					when "110111101001110" => rgb <= "101111";
					when "110111101001111" => rgb <= "101111";
					when "110111101010000" => rgb <= "101111";
					when "110111101010001" => rgb <= "101111";
					when "110111101010010" => rgb <= "101111";
					when "110111101010011" => rgb <= "101111";
					when "110111101010100" => rgb <= "101111";
					when "110111101010101" => rgb <= "101111";
					when "110111101010110" => rgb <= "101111";
					when "110111101010111" => rgb <= "101111";
					when "110111101011000" => rgb <= "101111";
					when "110111101011001" => rgb <= "101111";
					when "110111101011010" => rgb <= "101111";
					when "110111101011011" => rgb <= "101111";
					when "110111101011100" => rgb <= "101111";
					when "110111101011101" => rgb <= "101111";
					when "110111101011110" => rgb <= "101111";
					when "110111101011111" => rgb <= "101111";
					when "110111101100000" => rgb <= "101111";
					when "110111101100001" => rgb <= "101111";
					when "110111101100010" => rgb <= "101111";
					when "110111101100011" => rgb <= "101111";
					when "110111101100100" => rgb <= "101111";
					when "110111101100101" => rgb <= "101111";
					when "110111101100110" => rgb <= "101111";
					when "110111101100111" => rgb <= "101111";
					when "110111101101000" => rgb <= "101111";
					when "110111101101001" => rgb <= "101111";
					when "110111101101010" => rgb <= "101111";
					when "110111101101011" => rgb <= "101111";
					when "110111101101100" => rgb <= "101111";
					when "110111101101101" => rgb <= "101111";
					when "110111101101110" => rgb <= "101111";
					when "110111101101111" => rgb <= "101111";
					when "110111101110000" => rgb <= "101111";
					when "110111101110001" => rgb <= "101111";
					when "110111101110010" => rgb <= "101111";
					when "110111101110011" => rgb <= "101111";
					when "110111101110100" => rgb <= "101111";
					when "110111101110101" => rgb <= "101111";
					when "110111101110110" => rgb <= "101111";
					when "110111101110111" => rgb <= "101111";
					when "110111101111000" => rgb <= "101111";
					when "110111101111001" => rgb <= "101111";
					when "110111101111010" => rgb <= "101111";
					when "110111101111011" => rgb <= "101111";
					when "110111101111100" => rgb <= "101111";
					when "110111101111101" => rgb <= "101111";
					when "110111101111110" => rgb <= "101111";
					when "110111101111111" => rgb <= "101111";
					when "110111110000000" => rgb <= "101111";
					when "110111110000001" => rgb <= "101111";
					when "110111110000010" => rgb <= "101111";
					when "110111110000011" => rgb <= "101111";
					when "110111110000100" => rgb <= "101111";
					when "110111110000101" => rgb <= "101111";
					when "110111110000110" => rgb <= "101111";
					when "110111110000111" => rgb <= "101111";
					when "110111110001000" => rgb <= "101111";
					when "110111110001001" => rgb <= "101111";
					when "110111110001010" => rgb <= "101111";
					when "110111110001011" => rgb <= "101111";
					when "110111110001100" => rgb <= "101111";
					when "110111110001101" => rgb <= "101111";
					when "110111110001110" => rgb <= "101111";
					when "110111110001111" => rgb <= "101111";
					when "110111110010000" => rgb <= "101111";
					when "110111110010001" => rgb <= "101111";
					when "110111110010010" => rgb <= "101111";
					when "110111110010011" => rgb <= "101111";
					when "110111110010100" => rgb <= "101111";
					when "110111110010101" => rgb <= "101111";
					when "110111110010110" => rgb <= "101111";
					when "110111110010111" => rgb <= "101111";
					when "110111110011000" => rgb <= "101111";
					when "110111110011001" => rgb <= "101111";
					when "110111110011010" => rgb <= "101111";
					when "110111110011011" => rgb <= "101111";
					when "110111110011100" => rgb <= "101111";
					when "110111110011101" => rgb <= "101111";
					when "110111110011110" => rgb <= "101111";
					when "110111110011111" => rgb <= "101111";
					when "111000000000000" => rgb <= "101111";
					when "111000000000001" => rgb <= "101111";
					when "111000000000010" => rgb <= "101111";
					when "111000000000011" => rgb <= "101111";
					when "111000000000100" => rgb <= "101111";
					when "111000000000101" => rgb <= "101111";
					when "111000000000110" => rgb <= "101111";
					when "111000000000111" => rgb <= "101111";
					when "111000000001000" => rgb <= "101111";
					when "111000000001001" => rgb <= "101111";
					when "111000000001010" => rgb <= "101111";
					when "111000000001011" => rgb <= "101111";
					when "111000000001100" => rgb <= "101111";
					when "111000000001101" => rgb <= "101111";
					when "111000000001110" => rgb <= "101111";
					when "111000000001111" => rgb <= "101111";
					when "111000000010000" => rgb <= "101111";
					when "111000000010001" => rgb <= "101111";
					when "111000000010010" => rgb <= "101111";
					when "111000000010011" => rgb <= "101111";
					when "111000000010100" => rgb <= "101111";
					when "111000000010101" => rgb <= "101111";
					when "111000000010110" => rgb <= "101111";
					when "111000000010111" => rgb <= "101111";
					when "111000000011000" => rgb <= "000000";
					when "111000000011001" => rgb <= "000000";
					when "111000000011010" => rgb <= "000000";
					when "111000000011011" => rgb <= "000000";
					when "111000000011100" => rgb <= "100100";
					when "111000000011101" => rgb <= "100100";
					when "111000000011110" => rgb <= "100100";
					when "111000000011111" => rgb <= "100100";
					when "111000000100000" => rgb <= "100100";
					when "111000000100001" => rgb <= "100100";
					when "111000000100010" => rgb <= "100100";
					when "111000000100011" => rgb <= "100100";
					when "111000000100100" => rgb <= "100100";
					when "111000000100101" => rgb <= "100100";
					when "111000000100110" => rgb <= "100100";
					when "111000000100111" => rgb <= "100100";
					when "111000000101000" => rgb <= "100100";
					when "111000000101001" => rgb <= "100100";
					when "111000000101010" => rgb <= "100100";
					when "111000000101011" => rgb <= "100100";
					when "111000000101100" => rgb <= "100100";
					when "111000000101101" => rgb <= "100100";
					when "111000000101110" => rgb <= "100100";
					when "111000000101111" => rgb <= "100100";
					when "111000000110000" => rgb <= "100100";
					when "111000000110001" => rgb <= "100100";
					when "111000000110010" => rgb <= "100100";
					when "111000000110011" => rgb <= "100100";
					when "111000000110100" => rgb <= "100100";
					when "111000000110101" => rgb <= "100100";
					when "111000000110110" => rgb <= "100100";
					when "111000000110111" => rgb <= "100100";
					when "111000000111000" => rgb <= "100100";
					when "111000000111001" => rgb <= "100100";
					when "111000000111010" => rgb <= "010000";
					when "111000000111011" => rgb <= "010000";
					when "111000000111100" => rgb <= "000000";
					when "111000000111101" => rgb <= "000000";
					when "111000000111110" => rgb <= "000000";
					when "111000000111111" => rgb <= "000000";
					when "111000001000000" => rgb <= "101111";
					when "111000001000001" => rgb <= "101111";
					when "111000001000010" => rgb <= "101111";
					when "111000001000011" => rgb <= "101111";
					when "111000001000100" => rgb <= "101111";
					when "111000001000101" => rgb <= "101111";
					when "111000001000110" => rgb <= "101111";
					when "111000001000111" => rgb <= "101111";
					when "111000001001000" => rgb <= "101111";
					when "111000001001001" => rgb <= "101111";
					when "111000001001010" => rgb <= "101111";
					when "111000001001011" => rgb <= "101111";
					when "111000001001100" => rgb <= "101111";
					when "111000001001101" => rgb <= "101111";
					when "111000001001110" => rgb <= "101111";
					when "111000001001111" => rgb <= "101111";
					when "111000001010000" => rgb <= "101111";
					when "111000001010001" => rgb <= "101111";
					when "111000001010010" => rgb <= "101111";
					when "111000001010011" => rgb <= "101111";
					when "111000001010100" => rgb <= "101111";
					when "111000001010101" => rgb <= "101111";
					when "111000001010110" => rgb <= "101111";
					when "111000001010111" => rgb <= "101111";
					when "111000001011000" => rgb <= "101111";
					when "111000001011001" => rgb <= "101111";
					when "111000001011010" => rgb <= "101111";
					when "111000001011011" => rgb <= "101111";
					when "111000001011100" => rgb <= "101111";
					when "111000001011101" => rgb <= "101111";
					when "111000001011110" => rgb <= "101111";
					when "111000001011111" => rgb <= "101111";
					when "111000001100000" => rgb <= "101111";
					when "111000001100001" => rgb <= "101111";
					when "111000001100010" => rgb <= "101111";
					when "111000001100011" => rgb <= "101111";
					when "111000001100100" => rgb <= "101111";
					when "111000001100101" => rgb <= "101111";
					when "111000001100110" => rgb <= "101111";
					when "111000001100111" => rgb <= "101111";
					when "111000001101000" => rgb <= "101111";
					when "111000001101001" => rgb <= "101111";
					when "111000001101010" => rgb <= "101111";
					when "111000001101011" => rgb <= "101111";
					when "111000001101100" => rgb <= "101111";
					when "111000001101101" => rgb <= "101111";
					when "111000001101110" => rgb <= "101111";
					when "111000001101111" => rgb <= "101111";
					when "111000001110000" => rgb <= "101111";
					when "111000001110001" => rgb <= "101111";
					when "111000001110010" => rgb <= "101111";
					when "111000001110011" => rgb <= "101111";
					when "111000001110100" => rgb <= "101111";
					when "111000001110101" => rgb <= "101111";
					when "111000001110110" => rgb <= "101111";
					when "111000001110111" => rgb <= "101111";
					when "111000001111000" => rgb <= "101111";
					when "111000001111001" => rgb <= "101111";
					when "111000001111010" => rgb <= "101111";
					when "111000001111011" => rgb <= "101111";
					when "111000001111100" => rgb <= "101111";
					when "111000001111101" => rgb <= "101111";
					when "111000001111110" => rgb <= "101111";
					when "111000001111111" => rgb <= "101111";
					when "111000010000000" => rgb <= "101111";
					when "111000010000001" => rgb <= "101111";
					when "111000010000010" => rgb <= "101111";
					when "111000010000011" => rgb <= "101111";
					when "111000010000100" => rgb <= "101111";
					when "111000010000101" => rgb <= "101111";
					when "111000010000110" => rgb <= "101111";
					when "111000010000111" => rgb <= "101111";
					when "111000010001000" => rgb <= "101111";
					when "111000010001001" => rgb <= "101111";
					when "111000010001010" => rgb <= "101111";
					when "111000010001011" => rgb <= "101111";
					when "111000010001100" => rgb <= "101111";
					when "111000010001101" => rgb <= "101111";
					when "111000010001110" => rgb <= "101111";
					when "111000010001111" => rgb <= "101111";
					when "111000010010000" => rgb <= "101111";
					when "111000010010001" => rgb <= "101111";
					when "111000010010010" => rgb <= "101111";
					when "111000010010011" => rgb <= "101111";
					when "111000010010100" => rgb <= "101111";
					when "111000010010101" => rgb <= "101111";
					when "111000010010110" => rgb <= "101111";
					when "111000010010111" => rgb <= "101111";
					when "111000010011000" => rgb <= "101111";
					when "111000010011001" => rgb <= "101111";
					when "111000010011010" => rgb <= "101111";
					when "111000010011011" => rgb <= "101111";
					when "111000010011100" => rgb <= "101111";
					when "111000010011101" => rgb <= "101111";
					when "111000010011110" => rgb <= "101111";
					when "111000010011111" => rgb <= "101111";
					when "111000100000000" => rgb <= "101111";
					when "111000100000001" => rgb <= "101111";
					when "111000100000010" => rgb <= "101111";
					when "111000100000011" => rgb <= "101111";
					when "111000100000100" => rgb <= "101111";
					when "111000100000101" => rgb <= "101111";
					when "111000100000110" => rgb <= "101111";
					when "111000100000111" => rgb <= "101111";
					when "111000100001000" => rgb <= "101111";
					when "111000100001001" => rgb <= "101111";
					when "111000100001010" => rgb <= "101111";
					when "111000100001011" => rgb <= "101111";
					when "111000100001100" => rgb <= "101111";
					when "111000100001101" => rgb <= "101111";
					when "111000100001110" => rgb <= "101111";
					when "111000100001111" => rgb <= "101111";
					when "111000100010000" => rgb <= "101111";
					when "111000100010001" => rgb <= "101111";
					when "111000100010010" => rgb <= "101111";
					when "111000100010011" => rgb <= "101111";
					when "111000100010100" => rgb <= "101111";
					when "111000100010101" => rgb <= "101111";
					when "111000100010110" => rgb <= "101111";
					when "111000100010111" => rgb <= "101111";
					when "111000100011000" => rgb <= "000000";
					when "111000100011001" => rgb <= "000000";
					when "111000100011010" => rgb <= "000000";
					when "111000100011011" => rgb <= "000000";
					when "111000100011100" => rgb <= "100100";
					when "111000100011101" => rgb <= "100100";
					when "111000100011110" => rgb <= "100100";
					when "111000100011111" => rgb <= "100100";
					when "111000100100000" => rgb <= "100100";
					when "111000100100001" => rgb <= "100100";
					when "111000100100010" => rgb <= "100100";
					when "111000100100011" => rgb <= "100100";
					when "111000100100100" => rgb <= "100100";
					when "111000100100101" => rgb <= "100100";
					when "111000100100110" => rgb <= "100100";
					when "111000100100111" => rgb <= "100100";
					when "111000100101000" => rgb <= "100100";
					when "111000100101001" => rgb <= "100100";
					when "111000100101010" => rgb <= "100100";
					when "111000100101011" => rgb <= "100100";
					when "111000100101100" => rgb <= "100100";
					when "111000100101101" => rgb <= "100100";
					when "111000100101110" => rgb <= "100100";
					when "111000100101111" => rgb <= "100100";
					when "111000100110000" => rgb <= "100100";
					when "111000100110001" => rgb <= "100100";
					when "111000100110010" => rgb <= "100100";
					when "111000100110011" => rgb <= "100100";
					when "111000100110100" => rgb <= "100100";
					when "111000100110101" => rgb <= "100100";
					when "111000100110110" => rgb <= "100100";
					when "111000100110111" => rgb <= "100100";
					when "111000100111000" => rgb <= "100100";
					when "111000100111001" => rgb <= "100100";
					when "111000100111010" => rgb <= "010000";
					when "111000100111011" => rgb <= "010000";
					when "111000100111100" => rgb <= "000000";
					when "111000100111101" => rgb <= "000000";
					when "111000100111110" => rgb <= "000000";
					when "111000100111111" => rgb <= "000000";
					when "111000101000000" => rgb <= "101111";
					when "111000101000001" => rgb <= "101111";
					when "111000101000010" => rgb <= "101111";
					when "111000101000011" => rgb <= "101111";
					when "111000101000100" => rgb <= "101111";
					when "111000101000101" => rgb <= "101111";
					when "111000101000110" => rgb <= "101111";
					when "111000101000111" => rgb <= "101111";
					when "111000101001000" => rgb <= "101111";
					when "111000101001001" => rgb <= "101111";
					when "111000101001010" => rgb <= "101111";
					when "111000101001011" => rgb <= "101111";
					when "111000101001100" => rgb <= "101111";
					when "111000101001101" => rgb <= "101111";
					when "111000101001110" => rgb <= "101111";
					when "111000101001111" => rgb <= "101111";
					when "111000101010000" => rgb <= "101111";
					when "111000101010001" => rgb <= "101111";
					when "111000101010010" => rgb <= "101111";
					when "111000101010011" => rgb <= "101111";
					when "111000101010100" => rgb <= "101111";
					when "111000101010101" => rgb <= "101111";
					when "111000101010110" => rgb <= "101111";
					when "111000101010111" => rgb <= "101111";
					when "111000101011000" => rgb <= "101111";
					when "111000101011001" => rgb <= "101111";
					when "111000101011010" => rgb <= "101111";
					when "111000101011011" => rgb <= "101111";
					when "111000101011100" => rgb <= "101111";
					when "111000101011101" => rgb <= "101111";
					when "111000101011110" => rgb <= "101111";
					when "111000101011111" => rgb <= "101111";
					when "111000101100000" => rgb <= "101111";
					when "111000101100001" => rgb <= "101111";
					when "111000101100010" => rgb <= "101111";
					when "111000101100011" => rgb <= "101111";
					when "111000101100100" => rgb <= "101111";
					when "111000101100101" => rgb <= "101111";
					when "111000101100110" => rgb <= "101111";
					when "111000101100111" => rgb <= "101111";
					when "111000101101000" => rgb <= "101111";
					when "111000101101001" => rgb <= "101111";
					when "111000101101010" => rgb <= "101111";
					when "111000101101011" => rgb <= "101111";
					when "111000101101100" => rgb <= "101111";
					when "111000101101101" => rgb <= "101111";
					when "111000101101110" => rgb <= "101111";
					when "111000101101111" => rgb <= "101111";
					when "111000101110000" => rgb <= "101111";
					when "111000101110001" => rgb <= "101111";
					when "111000101110010" => rgb <= "101111";
					when "111000101110011" => rgb <= "101111";
					when "111000101110100" => rgb <= "101111";
					when "111000101110101" => rgb <= "101111";
					when "111000101110110" => rgb <= "101111";
					when "111000101110111" => rgb <= "101111";
					when "111000101111000" => rgb <= "101111";
					when "111000101111001" => rgb <= "101111";
					when "111000101111010" => rgb <= "101111";
					when "111000101111011" => rgb <= "101111";
					when "111000101111100" => rgb <= "101111";
					when "111000101111101" => rgb <= "101111";
					when "111000101111110" => rgb <= "101111";
					when "111000101111111" => rgb <= "101111";
					when "111000110000000" => rgb <= "101111";
					when "111000110000001" => rgb <= "101111";
					when "111000110000010" => rgb <= "101111";
					when "111000110000011" => rgb <= "101111";
					when "111000110000100" => rgb <= "101111";
					when "111000110000101" => rgb <= "101111";
					when "111000110000110" => rgb <= "101111";
					when "111000110000111" => rgb <= "101111";
					when "111000110001000" => rgb <= "101111";
					when "111000110001001" => rgb <= "101111";
					when "111000110001010" => rgb <= "101111";
					when "111000110001011" => rgb <= "101111";
					when "111000110001100" => rgb <= "101111";
					when "111000110001101" => rgb <= "101111";
					when "111000110001110" => rgb <= "101111";
					when "111000110001111" => rgb <= "101111";
					when "111000110010000" => rgb <= "101111";
					when "111000110010001" => rgb <= "101111";
					when "111000110010010" => rgb <= "101111";
					when "111000110010011" => rgb <= "101111";
					when "111000110010100" => rgb <= "101111";
					when "111000110010101" => rgb <= "101111";
					when "111000110010110" => rgb <= "101111";
					when "111000110010111" => rgb <= "101111";
					when "111000110011000" => rgb <= "101111";
					when "111000110011001" => rgb <= "101111";
					when "111000110011010" => rgb <= "101111";
					when "111000110011011" => rgb <= "101111";
					when "111000110011100" => rgb <= "101111";
					when "111000110011101" => rgb <= "101111";
					when "111000110011110" => rgb <= "101111";
					when "111000110011111" => rgb <= "101111";
					when "111001000000000" => rgb <= "101111";
					when "111001000000001" => rgb <= "101111";
					when "111001000000010" => rgb <= "101111";
					when "111001000000011" => rgb <= "101111";
					when "111001000000100" => rgb <= "101111";
					when "111001000000101" => rgb <= "101111";
					when "111001000000110" => rgb <= "101111";
					when "111001000000111" => rgb <= "101111";
					when "111001000001000" => rgb <= "101111";
					when "111001000001001" => rgb <= "101111";
					when "111001000001010" => rgb <= "101111";
					when "111001000001011" => rgb <= "101111";
					when "111001000001100" => rgb <= "101111";
					when "111001000001101" => rgb <= "101111";
					when "111001000001110" => rgb <= "101111";
					when "111001000001111" => rgb <= "101111";
					when "111001000010000" => rgb <= "101111";
					when "111001000010001" => rgb <= "101111";
					when "111001000010010" => rgb <= "000000";
					when "111001000010011" => rgb <= "000000";
					when "111001000010100" => rgb <= "000000";
					when "111001000010101" => rgb <= "000000";
					when "111001000010110" => rgb <= "000000";
					when "111001000010111" => rgb <= "000000";
					when "111001000011000" => rgb <= "000000";
					when "111001000011001" => rgb <= "000000";
					when "111001000011010" => rgb <= "000000";
					when "111001000011011" => rgb <= "000000";
					when "111001000011100" => rgb <= "000000";
					when "111001000011101" => rgb <= "000000";
					when "111001000011110" => rgb <= "000000";
					when "111001000011111" => rgb <= "000000";
					when "111001000100000" => rgb <= "000000";
					when "111001000100001" => rgb <= "000000";
					when "111001000100010" => rgb <= "000000";
					when "111001000100011" => rgb <= "000000";
					when "111001000100100" => rgb <= "000000";
					when "111001000100101" => rgb <= "000000";
					when "111001000100110" => rgb <= "000000";
					when "111001000100111" => rgb <= "000000";
					when "111001000101000" => rgb <= "000000";
					when "111001000101001" => rgb <= "000000";
					when "111001000101010" => rgb <= "000000";
					when "111001000101011" => rgb <= "000000";
					when "111001000101100" => rgb <= "000000";
					when "111001000101101" => rgb <= "000000";
					when "111001000101110" => rgb <= "000000";
					when "111001000101111" => rgb <= "000000";
					when "111001000110000" => rgb <= "000000";
					when "111001000110001" => rgb <= "000000";
					when "111001000110010" => rgb <= "000000";
					when "111001000110011" => rgb <= "000000";
					when "111001000110100" => rgb <= "000000";
					when "111001000110101" => rgb <= "000000";
					when "111001000110110" => rgb <= "000000";
					when "111001000110111" => rgb <= "000000";
					when "111001000111000" => rgb <= "000000";
					when "111001000111001" => rgb <= "000000";
					when "111001000111010" => rgb <= "000000";
					when "111001000111011" => rgb <= "000000";
					when "111001000111100" => rgb <= "000000";
					when "111001000111101" => rgb <= "000000";
					when "111001000111110" => rgb <= "000000";
					when "111001000111111" => rgb <= "000000";
					when "111001001000000" => rgb <= "000000";
					when "111001001000001" => rgb <= "000000";
					when "111001001000010" => rgb <= "000000";
					when "111001001000011" => rgb <= "000000";
					when "111001001000100" => rgb <= "000000";
					when "111001001000101" => rgb <= "000000";
					when "111001001000110" => rgb <= "101111";
					when "111001001000111" => rgb <= "101111";
					when "111001001001000" => rgb <= "101111";
					when "111001001001001" => rgb <= "101111";
					when "111001001001010" => rgb <= "101111";
					when "111001001001011" => rgb <= "101111";
					when "111001001001100" => rgb <= "101111";
					when "111001001001101" => rgb <= "101111";
					when "111001001001110" => rgb <= "101111";
					when "111001001001111" => rgb <= "101111";
					when "111001001010000" => rgb <= "101111";
					when "111001001010001" => rgb <= "101111";
					when "111001001010010" => rgb <= "101111";
					when "111001001010011" => rgb <= "101111";
					when "111001001010100" => rgb <= "101111";
					when "111001001010101" => rgb <= "101111";
					when "111001001010110" => rgb <= "101111";
					when "111001001010111" => rgb <= "101111";
					when "111001001011000" => rgb <= "101111";
					when "111001001011001" => rgb <= "101111";
					when "111001001011010" => rgb <= "101111";
					when "111001001011011" => rgb <= "101111";
					when "111001001011100" => rgb <= "101111";
					when "111001001011101" => rgb <= "101111";
					when "111001001011110" => rgb <= "101111";
					when "111001001011111" => rgb <= "101111";
					when "111001001100000" => rgb <= "101111";
					when "111001001100001" => rgb <= "101111";
					when "111001001100010" => rgb <= "101111";
					when "111001001100011" => rgb <= "101111";
					when "111001001100100" => rgb <= "101111";
					when "111001001100101" => rgb <= "101111";
					when "111001001100110" => rgb <= "101111";
					when "111001001100111" => rgb <= "101111";
					when "111001001101000" => rgb <= "101111";
					when "111001001101001" => rgb <= "101111";
					when "111001001101010" => rgb <= "101111";
					when "111001001101011" => rgb <= "101111";
					when "111001001101100" => rgb <= "101111";
					when "111001001101101" => rgb <= "101111";
					when "111001001101110" => rgb <= "101111";
					when "111001001101111" => rgb <= "101111";
					when "111001001110000" => rgb <= "101111";
					when "111001001110001" => rgb <= "101111";
					when "111001001110010" => rgb <= "101111";
					when "111001001110011" => rgb <= "101111";
					when "111001001110100" => rgb <= "101111";
					when "111001001110101" => rgb <= "101111";
					when "111001001110110" => rgb <= "101111";
					when "111001001110111" => rgb <= "101111";
					when "111001001111000" => rgb <= "101111";
					when "111001001111001" => rgb <= "101111";
					when "111001001111010" => rgb <= "101111";
					when "111001001111011" => rgb <= "101111";
					when "111001001111100" => rgb <= "101111";
					when "111001001111101" => rgb <= "101111";
					when "111001001111110" => rgb <= "101111";
					when "111001001111111" => rgb <= "101111";
					when "111001010000000" => rgb <= "101111";
					when "111001010000001" => rgb <= "101111";
					when "111001010000010" => rgb <= "101111";
					when "111001010000011" => rgb <= "101111";
					when "111001010000100" => rgb <= "101111";
					when "111001010000101" => rgb <= "101111";
					when "111001010000110" => rgb <= "101111";
					when "111001010000111" => rgb <= "101111";
					when "111001010001000" => rgb <= "101111";
					when "111001010001001" => rgb <= "101111";
					when "111001010001010" => rgb <= "101111";
					when "111001010001011" => rgb <= "101111";
					when "111001010001100" => rgb <= "101111";
					when "111001010001101" => rgb <= "101111";
					when "111001010001110" => rgb <= "101111";
					when "111001010001111" => rgb <= "101111";
					when "111001010010000" => rgb <= "101111";
					when "111001010010001" => rgb <= "101111";
					when "111001010010010" => rgb <= "101111";
					when "111001010010011" => rgb <= "101111";
					when "111001010010100" => rgb <= "101111";
					when "111001010010101" => rgb <= "101111";
					when "111001010010110" => rgb <= "101111";
					when "111001010010111" => rgb <= "101111";
					when "111001010011000" => rgb <= "101111";
					when "111001010011001" => rgb <= "101111";
					when "111001010011010" => rgb <= "101111";
					when "111001010011011" => rgb <= "101111";
					when "111001010011100" => rgb <= "101111";
					when "111001010011101" => rgb <= "101111";
					when "111001010011110" => rgb <= "101111";
					when "111001010011111" => rgb <= "101111";
					when "111001100000000" => rgb <= "101111";
					when "111001100000001" => rgb <= "101111";
					when "111001100000010" => rgb <= "101111";
					when "111001100000011" => rgb <= "101111";
					when "111001100000100" => rgb <= "101111";
					when "111001100000101" => rgb <= "101111";
					when "111001100000110" => rgb <= "101111";
					when "111001100000111" => rgb <= "101111";
					when "111001100001000" => rgb <= "101111";
					when "111001100001001" => rgb <= "101111";
					when "111001100001010" => rgb <= "101111";
					when "111001100001011" => rgb <= "101111";
					when "111001100001100" => rgb <= "101111";
					when "111001100001101" => rgb <= "101111";
					when "111001100001110" => rgb <= "101111";
					when "111001100001111" => rgb <= "101111";
					when "111001100010000" => rgb <= "101111";
					when "111001100010001" => rgb <= "101111";
					when "111001100010010" => rgb <= "000000";
					when "111001100010011" => rgb <= "000000";
					when "111001100010100" => rgb <= "000000";
					when "111001100010101" => rgb <= "000000";
					when "111001100010110" => rgb <= "000000";
					when "111001100010111" => rgb <= "000000";
					when "111001100011000" => rgb <= "000000";
					when "111001100011001" => rgb <= "000000";
					when "111001100011010" => rgb <= "000000";
					when "111001100011011" => rgb <= "000000";
					when "111001100011100" => rgb <= "000000";
					when "111001100011101" => rgb <= "000000";
					when "111001100011110" => rgb <= "000000";
					when "111001100011111" => rgb <= "000000";
					when "111001100100000" => rgb <= "000000";
					when "111001100100001" => rgb <= "000000";
					when "111001100100010" => rgb <= "000000";
					when "111001100100011" => rgb <= "000000";
					when "111001100100100" => rgb <= "000000";
					when "111001100100101" => rgb <= "000000";
					when "111001100100110" => rgb <= "000000";
					when "111001100100111" => rgb <= "000000";
					when "111001100101000" => rgb <= "000000";
					when "111001100101001" => rgb <= "000000";
					when "111001100101010" => rgb <= "000000";
					when "111001100101011" => rgb <= "000000";
					when "111001100101100" => rgb <= "000000";
					when "111001100101101" => rgb <= "000000";
					when "111001100101110" => rgb <= "000000";
					when "111001100101111" => rgb <= "000000";
					when "111001100110000" => rgb <= "000000";
					when "111001100110001" => rgb <= "000000";
					when "111001100110010" => rgb <= "000000";
					when "111001100110011" => rgb <= "000000";
					when "111001100110100" => rgb <= "000000";
					when "111001100110101" => rgb <= "000000";
					when "111001100110110" => rgb <= "000000";
					when "111001100110111" => rgb <= "000000";
					when "111001100111000" => rgb <= "000000";
					when "111001100111001" => rgb <= "000000";
					when "111001100111010" => rgb <= "000000";
					when "111001100111011" => rgb <= "000000";
					when "111001100111100" => rgb <= "000000";
					when "111001100111101" => rgb <= "000000";
					when "111001100111110" => rgb <= "000000";
					when "111001100111111" => rgb <= "000000";
					when "111001101000000" => rgb <= "000000";
					when "111001101000001" => rgb <= "000000";
					when "111001101000010" => rgb <= "000000";
					when "111001101000011" => rgb <= "000000";
					when "111001101000100" => rgb <= "000000";
					when "111001101000101" => rgb <= "000000";
					when "111001101000110" => rgb <= "101111";
					when "111001101000111" => rgb <= "101111";
					when "111001101001000" => rgb <= "101111";
					when "111001101001001" => rgb <= "101111";
					when "111001101001010" => rgb <= "101111";
					when "111001101001011" => rgb <= "101111";
					when "111001101001100" => rgb <= "101111";
					when "111001101001101" => rgb <= "101111";
					when "111001101001110" => rgb <= "101111";
					when "111001101001111" => rgb <= "101111";
					when "111001101010000" => rgb <= "101111";
					when "111001101010001" => rgb <= "101111";
					when "111001101010010" => rgb <= "101111";
					when "111001101010011" => rgb <= "101111";
					when "111001101010100" => rgb <= "101111";
					when "111001101010101" => rgb <= "101111";
					when "111001101010110" => rgb <= "101111";
					when "111001101010111" => rgb <= "101111";
					when "111001101011000" => rgb <= "101111";
					when "111001101011001" => rgb <= "101111";
					when "111001101011010" => rgb <= "101111";
					when "111001101011011" => rgb <= "101111";
					when "111001101011100" => rgb <= "101111";
					when "111001101011101" => rgb <= "101111";
					when "111001101011110" => rgb <= "101111";
					when "111001101011111" => rgb <= "101111";
					when "111001101100000" => rgb <= "101111";
					when "111001101100001" => rgb <= "101111";
					when "111001101100010" => rgb <= "101111";
					when "111001101100011" => rgb <= "101111";
					when "111001101100100" => rgb <= "101111";
					when "111001101100101" => rgb <= "101111";
					when "111001101100110" => rgb <= "101111";
					when "111001101100111" => rgb <= "101111";
					when "111001101101000" => rgb <= "101111";
					when "111001101101001" => rgb <= "101111";
					when "111001101101010" => rgb <= "101111";
					when "111001101101011" => rgb <= "101111";
					when "111001101101100" => rgb <= "101111";
					when "111001101101101" => rgb <= "101111";
					when "111001101101110" => rgb <= "101111";
					when "111001101101111" => rgb <= "101111";
					when "111001101110000" => rgb <= "101111";
					when "111001101110001" => rgb <= "101111";
					when "111001101110010" => rgb <= "101111";
					when "111001101110011" => rgb <= "101111";
					when "111001101110100" => rgb <= "101111";
					when "111001101110101" => rgb <= "101111";
					when "111001101110110" => rgb <= "101111";
					when "111001101110111" => rgb <= "101111";
					when "111001101111000" => rgb <= "101111";
					when "111001101111001" => rgb <= "101111";
					when "111001101111010" => rgb <= "101111";
					when "111001101111011" => rgb <= "101111";
					when "111001101111100" => rgb <= "101111";
					when "111001101111101" => rgb <= "101111";
					when "111001101111110" => rgb <= "101111";
					when "111001101111111" => rgb <= "101111";
					when "111001110000000" => rgb <= "101111";
					when "111001110000001" => rgb <= "101111";
					when "111001110000010" => rgb <= "101111";
					when "111001110000011" => rgb <= "101111";
					when "111001110000100" => rgb <= "101111";
					when "111001110000101" => rgb <= "101111";
					when "111001110000110" => rgb <= "101111";
					when "111001110000111" => rgb <= "101111";
					when "111001110001000" => rgb <= "101111";
					when "111001110001001" => rgb <= "101111";
					when "111001110001010" => rgb <= "101111";
					when "111001110001011" => rgb <= "101111";
					when "111001110001100" => rgb <= "101111";
					when "111001110001101" => rgb <= "101111";
					when "111001110001110" => rgb <= "101111";
					when "111001110001111" => rgb <= "101111";
					when "111001110010000" => rgb <= "101111";
					when "111001110010001" => rgb <= "101111";
					when "111001110010010" => rgb <= "101111";
					when "111001110010011" => rgb <= "101111";
					when "111001110010100" => rgb <= "101111";
					when "111001110010101" => rgb <= "101111";
					when "111001110010110" => rgb <= "101111";
					when "111001110010111" => rgb <= "101111";
					when "111001110011000" => rgb <= "101111";
					when "111001110011001" => rgb <= "101111";
					when "111001110011010" => rgb <= "101111";
					when "111001110011011" => rgb <= "101111";
					when "111001110011100" => rgb <= "101111";
					when "111001110011101" => rgb <= "101111";
					when "111001110011110" => rgb <= "101111";
					when "111001110011111" => rgb <= "101111";
					when "111010000000000" => rgb <= "011101";
					when "111010000000001" => rgb <= "011101";
					when "111010000000010" => rgb <= "001000";
					when "111010000000011" => rgb <= "001000";
					when "111010000000100" => rgb <= "101110";
					when "111010000000101" => rgb <= "101110";
					when "111010000000110" => rgb <= "011101";
					when "111010000000111" => rgb <= "011101";
					when "111010000001000" => rgb <= "101110";
					when "111010000001001" => rgb <= "101110";
					when "111010000001010" => rgb <= "001000";
					when "111010000001011" => rgb <= "001000";
					when "111010000001100" => rgb <= "011101";
					when "111010000001101" => rgb <= "011101";
					when "111010000001110" => rgb <= "001000";
					when "111010000001111" => rgb <= "001000";
					when "111010000010000" => rgb <= "011101";
					when "111010000010001" => rgb <= "011101";
					when "111010000010010" => rgb <= "000100";
					when "111010000010011" => rgb <= "000100";
					when "111010000010100" => rgb <= "011101";
					when "111010000010101" => rgb <= "011101";
					when "111010000010110" => rgb <= "011101";
					when "111010000010111" => rgb <= "011101";
					when "111010000011000" => rgb <= "101110";
					when "111010000011001" => rgb <= "101110";
					when "111010000011010" => rgb <= "011101";
					when "111010000011011" => rgb <= "011101";
					when "111010000011100" => rgb <= "011101";
					when "111010000011101" => rgb <= "011101";
					when "111010000011110" => rgb <= "011101";
					when "111010000011111" => rgb <= "011101";
					when "111010000100000" => rgb <= "011101";
					when "111010000100001" => rgb <= "011101";
					when "111010000100010" => rgb <= "001000";
					when "111010000100011" => rgb <= "001000";
					when "111010000100100" => rgb <= "000100";
					when "111010000100101" => rgb <= "000100";
					when "111010000100110" => rgb <= "011101";
					when "111010000100111" => rgb <= "011101";
					when "111010000101000" => rgb <= "011101";
					when "111010000101001" => rgb <= "011101";
					when "111010000101010" => rgb <= "000100";
					when "111010000101011" => rgb <= "000100";
					when "111010000101100" => rgb <= "011101";
					when "111010000101101" => rgb <= "011101";
					when "111010000101110" => rgb <= "011101";
					when "111010000101111" => rgb <= "011101";
					when "111010000110000" => rgb <= "011101";
					when "111010000110001" => rgb <= "011101";
					when "111010000110010" => rgb <= "101110";
					when "111010000110011" => rgb <= "101110";
					when "111010000110100" => rgb <= "011101";
					when "111010000110101" => rgb <= "011101";
					when "111010000110110" => rgb <= "011101";
					when "111010000110111" => rgb <= "011101";
					when "111010000111000" => rgb <= "011101";
					when "111010000111001" => rgb <= "011101";
					when "111010000111010" => rgb <= "001000";
					when "111010000111011" => rgb <= "001000";
					when "111010000111100" => rgb <= "011101";
					when "111010000111101" => rgb <= "011101";
					when "111010000111110" => rgb <= "101110";
					when "111010000111111" => rgb <= "101110";
					when "111010001000000" => rgb <= "011101";
					when "111010001000001" => rgb <= "011101";
					when "111010001000010" => rgb <= "011101";
					when "111010001000011" => rgb <= "011101";
					when "111010001000100" => rgb <= "000100";
					when "111010001000101" => rgb <= "000100";
					when "111010001000110" => rgb <= "011101";
					when "111010001000111" => rgb <= "011101";
					when "111010001001000" => rgb <= "001000";
					when "111010001001001" => rgb <= "001000";
					when "111010001001010" => rgb <= "011101";
					when "111010001001011" => rgb <= "011101";
					when "111010001001100" => rgb <= "101110";
					when "111010001001101" => rgb <= "101110";
					when "111010001001110" => rgb <= "011101";
					when "111010001001111" => rgb <= "011101";
					when "111010001010000" => rgb <= "011101";
					when "111010001010001" => rgb <= "011101";
					when "111010001010010" => rgb <= "011101";
					when "111010001010011" => rgb <= "011101";
					when "111010001010100" => rgb <= "000100";
					when "111010001010101" => rgb <= "000100";
					when "111010001010110" => rgb <= "011101";
					when "111010001010111" => rgb <= "011101";
					when "111010001011000" => rgb <= "011101";
					when "111010001011001" => rgb <= "011101";
					when "111010001011010" => rgb <= "001000";
					when "111010001011011" => rgb <= "001000";
					when "111010001011100" => rgb <= "011101";
					when "111010001011101" => rgb <= "011101";
					when "111010001011110" => rgb <= "101110";
					when "111010001011111" => rgb <= "101110";
					when "111010001100000" => rgb <= "011101";
					when "111010001100001" => rgb <= "011101";
					when "111010001100010" => rgb <= "001000";
					when "111010001100011" => rgb <= "001000";
					when "111010001100100" => rgb <= "011101";
					when "111010001100101" => rgb <= "011101";
					when "111010001100110" => rgb <= "101110";
					when "111010001100111" => rgb <= "101110";
					when "111010001101000" => rgb <= "011101";
					when "111010001101001" => rgb <= "011101";
					when "111010001101010" => rgb <= "101110";
					when "111010001101011" => rgb <= "101110";
					when "111010001101100" => rgb <= "101110";
					when "111010001101101" => rgb <= "101110";
					when "111010001101110" => rgb <= "011101";
					when "111010001101111" => rgb <= "011101";
					when "111010001110000" => rgb <= "001000";
					when "111010001110001" => rgb <= "001000";
					when "111010001110010" => rgb <= "011101";
					when "111010001110011" => rgb <= "011101";
					when "111010001110100" => rgb <= "000100";
					when "111010001110101" => rgb <= "000100";
					when "111010001110110" => rgb <= "001000";
					when "111010001110111" => rgb <= "001000";
					when "111010001111000" => rgb <= "011101";
					when "111010001111001" => rgb <= "011101";
					when "111010001111010" => rgb <= "011101";
					when "111010001111011" => rgb <= "011101";
					when "111010001111100" => rgb <= "000100";
					when "111010001111101" => rgb <= "000100";
					when "111010001111110" => rgb <= "011101";
					when "111010001111111" => rgb <= "011101";
					when "111010010000000" => rgb <= "101110";
					when "111010010000001" => rgb <= "101110";
					when "111010010000010" => rgb <= "011101";
					when "111010010000011" => rgb <= "011101";
					when "111010010000100" => rgb <= "011101";
					when "111010010000101" => rgb <= "011101";
					when "111010010000110" => rgb <= "001000";
					when "111010010000111" => rgb <= "001000";
					when "111010010001000" => rgb <= "011101";
					when "111010010001001" => rgb <= "011101";
					when "111010010001010" => rgb <= "101110";
					when "111010010001011" => rgb <= "101110";
					when "111010010001100" => rgb <= "011101";
					when "111010010001101" => rgb <= "011101";
					when "111010010001110" => rgb <= "011101";
					when "111010010001111" => rgb <= "011101";
					when "111010010010000" => rgb <= "000100";
					when "111010010010001" => rgb <= "000100";
					when "111010010010010" => rgb <= "011101";
					when "111010010010011" => rgb <= "011101";
					when "111010010010100" => rgb <= "001000";
					when "111010010010101" => rgb <= "001000";
					when "111010010010110" => rgb <= "011101";
					when "111010010010111" => rgb <= "011101";
					when "111010010011000" => rgb <= "101110";
					when "111010010011001" => rgb <= "101110";
					when "111010010011010" => rgb <= "011101";
					when "111010010011011" => rgb <= "011101";
					when "111010010011100" => rgb <= "001000";
					when "111010010011101" => rgb <= "001000";
					when "111010010011110" => rgb <= "011101";
					when "111010010011111" => rgb <= "011101";
					when "111010100000000" => rgb <= "011101";
					when "111010100000001" => rgb <= "011101";
					when "111010100000010" => rgb <= "001000";
					when "111010100000011" => rgb <= "001000";
					when "111010100000100" => rgb <= "101110";
					when "111010100000101" => rgb <= "101110";
					when "111010100000110" => rgb <= "011101";
					when "111010100000111" => rgb <= "011101";
					when "111010100001000" => rgb <= "101110";
					when "111010100001001" => rgb <= "101110";
					when "111010100001010" => rgb <= "001000";
					when "111010100001011" => rgb <= "001000";
					when "111010100001100" => rgb <= "011101";
					when "111010100001101" => rgb <= "011101";
					when "111010100001110" => rgb <= "001000";
					when "111010100001111" => rgb <= "001000";
					when "111010100010000" => rgb <= "011101";
					when "111010100010001" => rgb <= "011101";
					when "111010100010010" => rgb <= "000100";
					when "111010100010011" => rgb <= "000100";
					when "111010100010100" => rgb <= "011101";
					when "111010100010101" => rgb <= "011101";
					when "111010100010110" => rgb <= "011101";
					when "111010100010111" => rgb <= "011101";
					when "111010100011000" => rgb <= "101110";
					when "111010100011001" => rgb <= "101110";
					when "111010100011010" => rgb <= "011101";
					when "111010100011011" => rgb <= "011101";
					when "111010100011100" => rgb <= "011101";
					when "111010100011101" => rgb <= "011101";
					when "111010100011110" => rgb <= "011101";
					when "111010100011111" => rgb <= "011101";
					when "111010100100000" => rgb <= "011101";
					when "111010100100001" => rgb <= "011101";
					when "111010100100010" => rgb <= "001000";
					when "111010100100011" => rgb <= "001000";
					when "111010100100100" => rgb <= "000100";
					when "111010100100101" => rgb <= "000100";
					when "111010100100110" => rgb <= "011101";
					when "111010100100111" => rgb <= "011101";
					when "111010100101000" => rgb <= "011101";
					when "111010100101001" => rgb <= "011101";
					when "111010100101010" => rgb <= "000100";
					when "111010100101011" => rgb <= "000100";
					when "111010100101100" => rgb <= "011101";
					when "111010100101101" => rgb <= "011101";
					when "111010100101110" => rgb <= "011101";
					when "111010100101111" => rgb <= "011101";
					when "111010100110000" => rgb <= "011101";
					when "111010100110001" => rgb <= "011101";
					when "111010100110010" => rgb <= "101110";
					when "111010100110011" => rgb <= "101110";
					when "111010100110100" => rgb <= "011101";
					when "111010100110101" => rgb <= "011101";
					when "111010100110110" => rgb <= "011101";
					when "111010100110111" => rgb <= "011101";
					when "111010100111000" => rgb <= "011101";
					when "111010100111001" => rgb <= "011101";
					when "111010100111010" => rgb <= "001000";
					when "111010100111011" => rgb <= "001000";
					when "111010100111100" => rgb <= "011101";
					when "111010100111101" => rgb <= "011101";
					when "111010100111110" => rgb <= "101110";
					when "111010100111111" => rgb <= "101110";
					when "111010101000000" => rgb <= "011101";
					when "111010101000001" => rgb <= "011101";
					when "111010101000010" => rgb <= "011101";
					when "111010101000011" => rgb <= "011101";
					when "111010101000100" => rgb <= "000100";
					when "111010101000101" => rgb <= "000100";
					when "111010101000110" => rgb <= "011101";
					when "111010101000111" => rgb <= "011101";
					when "111010101001000" => rgb <= "001000";
					when "111010101001001" => rgb <= "001000";
					when "111010101001010" => rgb <= "011101";
					when "111010101001011" => rgb <= "011101";
					when "111010101001100" => rgb <= "101110";
					when "111010101001101" => rgb <= "101110";
					when "111010101001110" => rgb <= "011101";
					when "111010101001111" => rgb <= "011101";
					when "111010101010000" => rgb <= "011101";
					when "111010101010001" => rgb <= "011101";
					when "111010101010010" => rgb <= "011101";
					when "111010101010011" => rgb <= "011101";
					when "111010101010100" => rgb <= "000100";
					when "111010101010101" => rgb <= "000100";
					when "111010101010110" => rgb <= "011101";
					when "111010101010111" => rgb <= "011101";
					when "111010101011000" => rgb <= "011101";
					when "111010101011001" => rgb <= "011101";
					when "111010101011010" => rgb <= "001000";
					when "111010101011011" => rgb <= "001000";
					when "111010101011100" => rgb <= "011101";
					when "111010101011101" => rgb <= "011101";
					when "111010101011110" => rgb <= "101110";
					when "111010101011111" => rgb <= "101110";
					when "111010101100000" => rgb <= "011101";
					when "111010101100001" => rgb <= "011101";
					when "111010101100010" => rgb <= "001000";
					when "111010101100011" => rgb <= "001000";
					when "111010101100100" => rgb <= "011101";
					when "111010101100101" => rgb <= "011101";
					when "111010101100110" => rgb <= "101110";
					when "111010101100111" => rgb <= "101110";
					when "111010101101000" => rgb <= "011101";
					when "111010101101001" => rgb <= "011101";
					when "111010101101010" => rgb <= "101110";
					when "111010101101011" => rgb <= "101110";
					when "111010101101100" => rgb <= "101110";
					when "111010101101101" => rgb <= "101110";
					when "111010101101110" => rgb <= "011101";
					when "111010101101111" => rgb <= "011101";
					when "111010101110000" => rgb <= "001000";
					when "111010101110001" => rgb <= "001000";
					when "111010101110010" => rgb <= "011101";
					when "111010101110011" => rgb <= "011101";
					when "111010101110100" => rgb <= "000100";
					when "111010101110101" => rgb <= "000100";
					when "111010101110110" => rgb <= "001000";
					when "111010101110111" => rgb <= "001000";
					when "111010101111000" => rgb <= "011101";
					when "111010101111001" => rgb <= "011101";
					when "111010101111010" => rgb <= "011101";
					when "111010101111011" => rgb <= "011101";
					when "111010101111100" => rgb <= "000100";
					when "111010101111101" => rgb <= "000100";
					when "111010101111110" => rgb <= "011101";
					when "111010101111111" => rgb <= "011101";
					when "111010110000000" => rgb <= "101110";
					when "111010110000001" => rgb <= "101110";
					when "111010110000010" => rgb <= "011101";
					when "111010110000011" => rgb <= "011101";
					when "111010110000100" => rgb <= "011101";
					when "111010110000101" => rgb <= "011101";
					when "111010110000110" => rgb <= "001000";
					when "111010110000111" => rgb <= "001000";
					when "111010110001000" => rgb <= "011101";
					when "111010110001001" => rgb <= "011101";
					when "111010110001010" => rgb <= "101110";
					when "111010110001011" => rgb <= "101110";
					when "111010110001100" => rgb <= "011101";
					when "111010110001101" => rgb <= "011101";
					when "111010110001110" => rgb <= "011101";
					when "111010110001111" => rgb <= "011101";
					when "111010110010000" => rgb <= "000100";
					when "111010110010001" => rgb <= "000100";
					when "111010110010010" => rgb <= "011101";
					when "111010110010011" => rgb <= "011101";
					when "111010110010100" => rgb <= "001000";
					when "111010110010101" => rgb <= "001000";
					when "111010110010110" => rgb <= "011101";
					when "111010110010111" => rgb <= "011101";
					when "111010110011000" => rgb <= "101110";
					when "111010110011001" => rgb <= "101110";
					when "111010110011010" => rgb <= "011101";
					when "111010110011011" => rgb <= "011101";
					when "111010110011100" => rgb <= "001000";
					when "111010110011101" => rgb <= "001000";
					when "111010110011110" => rgb <= "011101";
					when "111010110011111" => rgb <= "011101";
					when "111011000000000" => rgb <= "011101";
					when "111011000000001" => rgb <= "011101";
					when "111011000000010" => rgb <= "011101";
					when "111011000000011" => rgb <= "011101";
					when "111011000000100" => rgb <= "001000";
					when "111011000000101" => rgb <= "001000";
					when "111011000000110" => rgb <= "011101";
					when "111011000000111" => rgb <= "011101";
					when "111011000001000" => rgb <= "000100";
					when "111011000001001" => rgb <= "000100";
					when "111011000001010" => rgb <= "011101";
					when "111011000001011" => rgb <= "011101";
					when "111011000001100" => rgb <= "101110";
					when "111011000001101" => rgb <= "101110";
					when "111011000001110" => rgb <= "011101";
					when "111011000001111" => rgb <= "011101";
					when "111011000010000" => rgb <= "011101";
					when "111011000010001" => rgb <= "011101";
					when "111011000010010" => rgb <= "011101";
					when "111011000010011" => rgb <= "011101";
					when "111011000010100" => rgb <= "011101";
					when "111011000010101" => rgb <= "011101";
					when "111011000010110" => rgb <= "001000";
					when "111011000010111" => rgb <= "001000";
					when "111011000011000" => rgb <= "011101";
					when "111011000011001" => rgb <= "011101";
					when "111011000011010" => rgb <= "000100";
					when "111011000011011" => rgb <= "000100";
					when "111011000011100" => rgb <= "011101";
					when "111011000011101" => rgb <= "011101";
					when "111011000011110" => rgb <= "011101";
					when "111011000011111" => rgb <= "011101";
					when "111011000100000" => rgb <= "001000";
					when "111011000100001" => rgb <= "001000";
					when "111011000100010" => rgb <= "011101";
					when "111011000100011" => rgb <= "011101";
					when "111011000100100" => rgb <= "101110";
					when "111011000100101" => rgb <= "101110";
					when "111011000100110" => rgb <= "101110";
					when "111011000100111" => rgb <= "101110";
					when "111011000101000" => rgb <= "101110";
					when "111011000101001" => rgb <= "101110";
					when "111011000101010" => rgb <= "011101";
					when "111011000101011" => rgb <= "011101";
					when "111011000101100" => rgb <= "011101";
					when "111011000101101" => rgb <= "011101";
					when "111011000101110" => rgb <= "011101";
					when "111011000101111" => rgb <= "011101";
					when "111011000110000" => rgb <= "000100";
					when "111011000110001" => rgb <= "000100";
					when "111011000110010" => rgb <= "000100";
					when "111011000110011" => rgb <= "000100";
					when "111011000110100" => rgb <= "011101";
					when "111011000110101" => rgb <= "011101";
					when "111011000110110" => rgb <= "001000";
					when "111011000110111" => rgb <= "001000";
					when "111011000111000" => rgb <= "001000";
					when "111011000111001" => rgb <= "001000";
					when "111011000111010" => rgb <= "011101";
					when "111011000111011" => rgb <= "011101";
					when "111011000111100" => rgb <= "011101";
					when "111011000111101" => rgb <= "011101";
					when "111011000111110" => rgb <= "011101";
					when "111011000111111" => rgb <= "011101";
					when "111011001000000" => rgb <= "011101";
					when "111011001000001" => rgb <= "011101";
					when "111011001000010" => rgb <= "101110";
					when "111011001000011" => rgb <= "101110";
					when "111011001000100" => rgb <= "011101";
					when "111011001000101" => rgb <= "011101";
					when "111011001000110" => rgb <= "011101";
					when "111011001000111" => rgb <= "011101";
					when "111011001001000" => rgb <= "000100";
					when "111011001001001" => rgb <= "000100";
					when "111011001001010" => rgb <= "011101";
					when "111011001001011" => rgb <= "011101";
					when "111011001001100" => rgb <= "011101";
					when "111011001001101" => rgb <= "011101";
					when "111011001001110" => rgb <= "011101";
					when "111011001001111" => rgb <= "011101";
					when "111011001010000" => rgb <= "000100";
					when "111011001010001" => rgb <= "000100";
					when "111011001010010" => rgb <= "011101";
					when "111011001010011" => rgb <= "011101";
					when "111011001010100" => rgb <= "101110";
					when "111011001010101" => rgb <= "101110";
					when "111011001010110" => rgb <= "011101";
					when "111011001010111" => rgb <= "011101";
					when "111011001011000" => rgb <= "011101";
					when "111011001011001" => rgb <= "011101";
					when "111011001011010" => rgb <= "011101";
					when "111011001011011" => rgb <= "011101";
					when "111011001011100" => rgb <= "000100";
					when "111011001011101" => rgb <= "000100";
					when "111011001011110" => rgb <= "011101";
					when "111011001011111" => rgb <= "011101";
					when "111011001100000" => rgb <= "001000";
					when "111011001100001" => rgb <= "001000";
					when "111011001100010" => rgb <= "011101";
					when "111011001100011" => rgb <= "011101";
					when "111011001100100" => rgb <= "011101";
					when "111011001100101" => rgb <= "011101";
					when "111011001100110" => rgb <= "011101";
					when "111011001100111" => rgb <= "011101";
					when "111011001101000" => rgb <= "000100";
					when "111011001101001" => rgb <= "000100";
					when "111011001101010" => rgb <= "011101";
					when "111011001101011" => rgb <= "011101";
					when "111011001101100" => rgb <= "101110";
					when "111011001101101" => rgb <= "101110";
					when "111011001101110" => rgb <= "011101";
					when "111011001101111" => rgb <= "011101";
					when "111011001110000" => rgb <= "011101";
					when "111011001110001" => rgb <= "011101";
					when "111011001110010" => rgb <= "000100";
					when "111011001110011" => rgb <= "000100";
					when "111011001110100" => rgb <= "000100";
					when "111011001110101" => rgb <= "000100";
					when "111011001110110" => rgb <= "011101";
					when "111011001110111" => rgb <= "011101";
					when "111011001111000" => rgb <= "101110";
					when "111011001111001" => rgb <= "101110";
					when "111011001111010" => rgb <= "011101";
					when "111011001111011" => rgb <= "011101";
					when "111011001111100" => rgb <= "001000";
					when "111011001111101" => rgb <= "001000";
					when "111011001111110" => rgb <= "011101";
					when "111011001111111" => rgb <= "011101";
					when "111011010000000" => rgb <= "011101";
					when "111011010000001" => rgb <= "011101";
					when "111011010000010" => rgb <= "011101";
					when "111011010000011" => rgb <= "011101";
					when "111011010000100" => rgb <= "101110";
					when "111011010000101" => rgb <= "101110";
					when "111011010000110" => rgb <= "001000";
					when "111011010000111" => rgb <= "001000";
					when "111011010001000" => rgb <= "001000";
					when "111011010001001" => rgb <= "001000";
					when "111011010001010" => rgb <= "011101";
					when "111011010001011" => rgb <= "011101";
					when "111011010001100" => rgb <= "101110";
					when "111011010001101" => rgb <= "101110";
					when "111011010001110" => rgb <= "011101";
					when "111011010001111" => rgb <= "011101";
					when "111011010010000" => rgb <= "000100";
					when "111011010010001" => rgb <= "000100";
					when "111011010010010" => rgb <= "011101";
					when "111011010010011" => rgb <= "011101";
					when "111011010010100" => rgb <= "011101";
					when "111011010010101" => rgb <= "011101";
					when "111011010010110" => rgb <= "101110";
					when "111011010010111" => rgb <= "101110";
					when "111011010011000" => rgb <= "001000";
					when "111011010011001" => rgb <= "001000";
					when "111011010011010" => rgb <= "011101";
					when "111011010011011" => rgb <= "011101";
					when "111011010011100" => rgb <= "000100";
					when "111011010011101" => rgb <= "000100";
					when "111011010011110" => rgb <= "011101";
					when "111011010011111" => rgb <= "011101";
					when "111011100000000" => rgb <= "011101";
					when "111011100000001" => rgb <= "011101";
					when "111011100000010" => rgb <= "011101";
					when "111011100000011" => rgb <= "011101";
					when "111011100000100" => rgb <= "001000";
					when "111011100000101" => rgb <= "001000";
					when "111011100000110" => rgb <= "011101";
					when "111011100000111" => rgb <= "011101";
					when "111011100001000" => rgb <= "000100";
					when "111011100001001" => rgb <= "000100";
					when "111011100001010" => rgb <= "011101";
					when "111011100001011" => rgb <= "011101";
					when "111011100001100" => rgb <= "101110";
					when "111011100001101" => rgb <= "101110";
					when "111011100001110" => rgb <= "011101";
					when "111011100001111" => rgb <= "011101";
					when "111011100010000" => rgb <= "011101";
					when "111011100010001" => rgb <= "011101";
					when "111011100010010" => rgb <= "011101";
					when "111011100010011" => rgb <= "011101";
					when "111011100010100" => rgb <= "011101";
					when "111011100010101" => rgb <= "011101";
					when "111011100010110" => rgb <= "001000";
					when "111011100010111" => rgb <= "001000";
					when "111011100011000" => rgb <= "011101";
					when "111011100011001" => rgb <= "011101";
					when "111011100011010" => rgb <= "000100";
					when "111011100011011" => rgb <= "000100";
					when "111011100011100" => rgb <= "011101";
					when "111011100011101" => rgb <= "011101";
					when "111011100011110" => rgb <= "011101";
					when "111011100011111" => rgb <= "011101";
					when "111011100100000" => rgb <= "001000";
					when "111011100100001" => rgb <= "001000";
					when "111011100100010" => rgb <= "011101";
					when "111011100100011" => rgb <= "011101";
					when "111011100100100" => rgb <= "101110";
					when "111011100100101" => rgb <= "101110";
					when "111011100100110" => rgb <= "101110";
					when "111011100100111" => rgb <= "101110";
					when "111011100101000" => rgb <= "101110";
					when "111011100101001" => rgb <= "101110";
					when "111011100101010" => rgb <= "011101";
					when "111011100101011" => rgb <= "011101";
					when "111011100101100" => rgb <= "011101";
					when "111011100101101" => rgb <= "011101";
					when "111011100101110" => rgb <= "011101";
					when "111011100101111" => rgb <= "011101";
					when "111011100110000" => rgb <= "000100";
					when "111011100110001" => rgb <= "000100";
					when "111011100110010" => rgb <= "000100";
					when "111011100110011" => rgb <= "000100";
					when "111011100110100" => rgb <= "011101";
					when "111011100110101" => rgb <= "011101";
					when "111011100110110" => rgb <= "001000";
					when "111011100110111" => rgb <= "001000";
					when "111011100111000" => rgb <= "001000";
					when "111011100111001" => rgb <= "001000";
					when "111011100111010" => rgb <= "011101";
					when "111011100111011" => rgb <= "011101";
					when "111011100111100" => rgb <= "011101";
					when "111011100111101" => rgb <= "011101";
					when "111011100111110" => rgb <= "011101";
					when "111011100111111" => rgb <= "011101";
					when "111011101000000" => rgb <= "011101";
					when "111011101000001" => rgb <= "011101";
					when "111011101000010" => rgb <= "101110";
					when "111011101000011" => rgb <= "101110";
					when "111011101000100" => rgb <= "011101";
					when "111011101000101" => rgb <= "011101";
					when "111011101000110" => rgb <= "011101";
					when "111011101000111" => rgb <= "011101";
					when "111011101001000" => rgb <= "000100";
					when "111011101001001" => rgb <= "000100";
					when "111011101001010" => rgb <= "011101";
					when "111011101001011" => rgb <= "011101";
					when "111011101001100" => rgb <= "011101";
					when "111011101001101" => rgb <= "011101";
					when "111011101001110" => rgb <= "011101";
					when "111011101001111" => rgb <= "011101";
					when "111011101010000" => rgb <= "000100";
					when "111011101010001" => rgb <= "000100";
					when "111011101010010" => rgb <= "011101";
					when "111011101010011" => rgb <= "011101";
					when "111011101010100" => rgb <= "101110";
					when "111011101010101" => rgb <= "101110";
					when "111011101010110" => rgb <= "011101";
					when "111011101010111" => rgb <= "011101";
					when "111011101011000" => rgb <= "011101";
					when "111011101011001" => rgb <= "011101";
					when "111011101011010" => rgb <= "011101";
					when "111011101011011" => rgb <= "011101";
					when "111011101011100" => rgb <= "000100";
					when "111011101011101" => rgb <= "000100";
					when "111011101011110" => rgb <= "011101";
					when "111011101011111" => rgb <= "011101";
					when "111011101100000" => rgb <= "001000";
					when "111011101100001" => rgb <= "001000";
					when "111011101100010" => rgb <= "011101";
					when "111011101100011" => rgb <= "011101";
					when "111011101100100" => rgb <= "011101";
					when "111011101100101" => rgb <= "011101";
					when "111011101100110" => rgb <= "011101";
					when "111011101100111" => rgb <= "011101";
					when "111011101101000" => rgb <= "000100";
					when "111011101101001" => rgb <= "000100";
					when "111011101101010" => rgb <= "011101";
					when "111011101101011" => rgb <= "011101";
					when "111011101101100" => rgb <= "101110";
					when "111011101101101" => rgb <= "101110";
					when "111011101101110" => rgb <= "011101";
					when "111011101101111" => rgb <= "011101";
					when "111011101110000" => rgb <= "011101";
					when "111011101110001" => rgb <= "011101";
					when "111011101110010" => rgb <= "000100";
					when "111011101110011" => rgb <= "000100";
					when "111011101110100" => rgb <= "000100";
					when "111011101110101" => rgb <= "000100";
					when "111011101110110" => rgb <= "011101";
					when "111011101110111" => rgb <= "011101";
					when "111011101111000" => rgb <= "101110";
					when "111011101111001" => rgb <= "101110";
					when "111011101111010" => rgb <= "011101";
					when "111011101111011" => rgb <= "011101";
					when "111011101111100" => rgb <= "001000";
					when "111011101111101" => rgb <= "001000";
					when "111011101111110" => rgb <= "011101";
					when "111011101111111" => rgb <= "011101";
					when "111011110000000" => rgb <= "011101";
					when "111011110000001" => rgb <= "011101";
					when "111011110000010" => rgb <= "011101";
					when "111011110000011" => rgb <= "011101";
					when "111011110000100" => rgb <= "101110";
					when "111011110000101" => rgb <= "101110";
					when "111011110000110" => rgb <= "001000";
					when "111011110000111" => rgb <= "001000";
					when "111011110001000" => rgb <= "001000";
					when "111011110001001" => rgb <= "001000";
					when "111011110001010" => rgb <= "011101";
					when "111011110001011" => rgb <= "011101";
					when "111011110001100" => rgb <= "101110";
					when "111011110001101" => rgb <= "101110";
					when "111011110001110" => rgb <= "011101";
					when "111011110001111" => rgb <= "011101";
					when "111011110010000" => rgb <= "000100";
					when "111011110010001" => rgb <= "000100";
					when "111011110010010" => rgb <= "011101";
					when "111011110010011" => rgb <= "011101";
					when "111011110010100" => rgb <= "011101";
					when "111011110010101" => rgb <= "011101";
					when "111011110010110" => rgb <= "101110";
					when "111011110010111" => rgb <= "101110";
					when "111011110011000" => rgb <= "001000";
					when "111011110011001" => rgb <= "001000";
					when "111011110011010" => rgb <= "011101";
					when "111011110011011" => rgb <= "011101";
					when "111011110011100" => rgb <= "000100";
					when "111011110011101" => rgb <= "000100";
					when "111011110011110" => rgb <= "011101";
					when "111011110011111" => rgb <= "011101";
					when others => rgb <= "000000";
		end case;
	end if;
   end process;
   totaladr <= std_logic_vector(yadr) & std_logic_vector(xadr);
end;