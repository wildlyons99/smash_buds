library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tony_run_rom2 is
  port(
	  clk : in std_logic;
	  xadr: in unsigned(4 downto 0);
	  yadr : in unsigned(5 downto 0); -- 0-1023
	  rgb : out std_logic_vector(5 downto 0)
      );
end tony_run_rom2;

architecture synth of tony_run_rom2 is
signal totaladr : std_logic_vector(10 downto 0);
begin
   process (clk) begin
	if rising_edge(clk) then
		case totaladr is
					when "00000000000" => rgb <= "110110";
					when "00000000001" => rgb <= "110110";
					when "00000000010" => rgb <= "110110";
					when "00000000011" => rgb <= "110110";
					when "00000000100" => rgb <= "110110";
					when "00000000101" => rgb <= "110110";
					when "00000000110" => rgb <= "110110";
					when "00000000111" => rgb <= "110110";
					when "00000001000" => rgb <= "110110";
					when "00000001001" => rgb <= "110110";
					when "00000001010" => rgb <= "110110";
					when "00000001011" => rgb <= "110110";
					when "00000001100" => rgb <= "110110";
					when "00000001101" => rgb <= "110110";
					when "00000001110" => rgb <= "110110";
					when "00000001111" => rgb <= "110110";
					when "00000010000" => rgb <= "110110";
					when "00000010001" => rgb <= "110110";
					when "00000010010" => rgb <= "110110";
					when "00000010011" => rgb <= "110110";
					when "00000010100" => rgb <= "110110";
					when "00000010101" => rgb <= "110110";
					when "00000010110" => rgb <= "110110";
					when "00000010111" => rgb <= "110110";
					when "00000011000" => rgb <= "110110";
					when "00000011001" => rgb <= "110110";
					when "00000100000" => rgb <= "110110";
					when "00000100001" => rgb <= "110110";
					when "00000100010" => rgb <= "110110";
					when "00000100011" => rgb <= "110110";
					when "00000100100" => rgb <= "110110";
					when "00000100101" => rgb <= "110110";
					when "00000100110" => rgb <= "110110";
					when "00000100111" => rgb <= "110110";
					when "00000101000" => rgb <= "110110";
					when "00000101001" => rgb <= "110110";
					when "00000101010" => rgb <= "110110";
					when "00000101011" => rgb <= "110110";
					when "00000101100" => rgb <= "110110";
					when "00000101101" => rgb <= "110110";
					when "00000101110" => rgb <= "110110";
					when "00000101111" => rgb <= "110110";
					when "00000110000" => rgb <= "110110";
					when "00000110001" => rgb <= "110110";
					when "00000110010" => rgb <= "110110";
					when "00000110011" => rgb <= "110110";
					when "00000110100" => rgb <= "110110";
					when "00000110101" => rgb <= "110110";
					when "00000110110" => rgb <= "110110";
					when "00000110111" => rgb <= "110110";
					when "00000111000" => rgb <= "110110";
					when "00000111001" => rgb <= "110110";
					when "00001000000" => rgb <= "110110";
					when "00001000001" => rgb <= "110110";
					when "00001000010" => rgb <= "110110";
					when "00001000011" => rgb <= "110110";
					when "00001000100" => rgb <= "101010";
					when "00001000101" => rgb <= "101010";
					when "00001000110" => rgb <= "101010";
					when "00001000111" => rgb <= "101010";
					when "00001001000" => rgb <= "101010";
					when "00001001001" => rgb <= "101010";
					when "00001001010" => rgb <= "101010";
					when "00001001011" => rgb <= "101010";
					when "00001001100" => rgb <= "101010";
					when "00001001101" => rgb <= "101010";
					when "00001001110" => rgb <= "101010";
					when "00001001111" => rgb <= "101010";
					when "00001010000" => rgb <= "101010";
					when "00001010001" => rgb <= "101010";
					when "00001010010" => rgb <= "101010";
					when "00001010011" => rgb <= "101010";
					when "00001010100" => rgb <= "101010";
					when "00001010101" => rgb <= "101010";
					when "00001010110" => rgb <= "110110";
					when "00001010111" => rgb <= "110110";
					when "00001011000" => rgb <= "110110";
					when "00001011001" => rgb <= "110110";
					when "00001100000" => rgb <= "110110";
					when "00001100001" => rgb <= "110110";
					when "00001100010" => rgb <= "110110";
					when "00001100011" => rgb <= "110110";
					when "00001100100" => rgb <= "101010";
					when "00001100101" => rgb <= "101010";
					when "00001100110" => rgb <= "101010";
					when "00001100111" => rgb <= "101010";
					when "00001101000" => rgb <= "101010";
					when "00001101001" => rgb <= "101010";
					when "00001101010" => rgb <= "101010";
					when "00001101011" => rgb <= "101010";
					when "00001101100" => rgb <= "101010";
					when "00001101101" => rgb <= "101010";
					when "00001101110" => rgb <= "101010";
					when "00001101111" => rgb <= "101010";
					when "00001110000" => rgb <= "101010";
					when "00001110001" => rgb <= "101010";
					when "00001110010" => rgb <= "101010";
					when "00001110011" => rgb <= "101010";
					when "00001110100" => rgb <= "101010";
					when "00001110101" => rgb <= "101010";
					when "00001110110" => rgb <= "110110";
					when "00001110111" => rgb <= "110110";
					when "00001111000" => rgb <= "110110";
					when "00001111001" => rgb <= "110110";
					when "00010000000" => rgb <= "110110";
					when "00010000001" => rgb <= "110110";
					when "00010000010" => rgb <= "101010";
					when "00010000011" => rgb <= "101010";
					when "00010000100" => rgb <= "101010";
					when "00010000101" => rgb <= "101010";
					when "00010000110" => rgb <= "101010";
					when "00010000111" => rgb <= "101010";
					when "00010001000" => rgb <= "101010";
					when "00010001001" => rgb <= "101010";
					when "00010001010" => rgb <= "101010";
					when "00010001011" => rgb <= "101010";
					when "00010001100" => rgb <= "101010";
					when "00010001101" => rgb <= "101010";
					when "00010001110" => rgb <= "101010";
					when "00010001111" => rgb <= "101010";
					when "00010010000" => rgb <= "101010";
					when "00010010001" => rgb <= "101010";
					when "00010010010" => rgb <= "101010";
					when "00010010011" => rgb <= "101010";
					when "00010010100" => rgb <= "101010";
					when "00010010101" => rgb <= "101010";
					when "00010010110" => rgb <= "101010";
					when "00010010111" => rgb <= "101010";
					when "00010011000" => rgb <= "110110";
					when "00010011001" => rgb <= "110110";
					when "00010100000" => rgb <= "110110";
					when "00010100001" => rgb <= "110110";
					when "00010100010" => rgb <= "101010";
					when "00010100011" => rgb <= "101010";
					when "00010100100" => rgb <= "101010";
					when "00010100101" => rgb <= "101010";
					when "00010100110" => rgb <= "101010";
					when "00010100111" => rgb <= "101010";
					when "00010101000" => rgb <= "101010";
					when "00010101001" => rgb <= "101010";
					when "00010101010" => rgb <= "101010";
					when "00010101011" => rgb <= "101010";
					when "00010101100" => rgb <= "101010";
					when "00010101101" => rgb <= "101010";
					when "00010101110" => rgb <= "101010";
					when "00010101111" => rgb <= "101010";
					when "00010110000" => rgb <= "101010";
					when "00010110001" => rgb <= "101010";
					when "00010110010" => rgb <= "101010";
					when "00010110011" => rgb <= "101010";
					when "00010110100" => rgb <= "101010";
					when "00010110101" => rgb <= "101010";
					when "00010110110" => rgb <= "101010";
					when "00010110111" => rgb <= "101010";
					when "00010111000" => rgb <= "110110";
					when "00010111001" => rgb <= "110110";
					when "00011000000" => rgb <= "101010";
					when "00011000001" => rgb <= "101010";
					when "00011000010" => rgb <= "101010";
					when "00011000011" => rgb <= "101010";
					when "00011000100" => rgb <= "101010";
					when "00011000101" => rgb <= "101010";
					when "00011000110" => rgb <= "101010";
					when "00011000111" => rgb <= "101010";
					when "00011001000" => rgb <= "111110";
					when "00011001001" => rgb <= "111110";
					when "00011001010" => rgb <= "111110";
					when "00011001011" => rgb <= "111110";
					when "00011001100" => rgb <= "111110";
					when "00011001101" => rgb <= "111110";
					when "00011001110" => rgb <= "111110";
					when "00011001111" => rgb <= "111110";
					when "00011010000" => rgb <= "111110";
					when "00011010001" => rgb <= "111110";
					when "00011010010" => rgb <= "101010";
					when "00011010011" => rgb <= "101010";
					when "00011010100" => rgb <= "101010";
					when "00011010101" => rgb <= "101010";
					when "00011010110" => rgb <= "101010";
					when "00011010111" => rgb <= "101010";
					when "00011011000" => rgb <= "110110";
					when "00011011001" => rgb <= "110110";
					when "00011100000" => rgb <= "101010";
					when "00011100001" => rgb <= "101010";
					when "00011100010" => rgb <= "101010";
					when "00011100011" => rgb <= "101010";
					when "00011100100" => rgb <= "101010";
					when "00011100101" => rgb <= "101010";
					when "00011100110" => rgb <= "101010";
					when "00011100111" => rgb <= "101010";
					when "00011101000" => rgb <= "111110";
					when "00011101001" => rgb <= "111110";
					when "00011101010" => rgb <= "111110";
					when "00011101011" => rgb <= "111110";
					when "00011101100" => rgb <= "111110";
					when "00011101101" => rgb <= "111110";
					when "00011101110" => rgb <= "111110";
					when "00011101111" => rgb <= "111110";
					when "00011110000" => rgb <= "111110";
					when "00011110001" => rgb <= "111110";
					when "00011110010" => rgb <= "101010";
					when "00011110011" => rgb <= "101010";
					when "00011110100" => rgb <= "101010";
					when "00011110101" => rgb <= "101010";
					when "00011110110" => rgb <= "101010";
					when "00011110111" => rgb <= "101010";
					when "00011111000" => rgb <= "110110";
					when "00011111001" => rgb <= "110110";
					when "00100000000" => rgb <= "101010";
					when "00100000001" => rgb <= "101010";
					when "00100000010" => rgb <= "101010";
					when "00100000011" => rgb <= "101010";
					when "00100000100" => rgb <= "101010";
					when "00100000101" => rgb <= "101010";
					when "00100000110" => rgb <= "111110";
					when "00100000111" => rgb <= "111110";
					when "00100001000" => rgb <= "111110";
					when "00100001001" => rgb <= "111110";
					when "00100001010" => rgb <= "111110";
					when "00100001011" => rgb <= "111110";
					when "00100001100" => rgb <= "111110";
					when "00100001101" => rgb <= "111110";
					when "00100001110" => rgb <= "111110";
					when "00100001111" => rgb <= "111110";
					when "00100010000" => rgb <= "111110";
					when "00100010001" => rgb <= "111110";
					when "00100010010" => rgb <= "111110";
					when "00100010011" => rgb <= "111110";
					when "00100010100" => rgb <= "111110";
					when "00100010101" => rgb <= "111110";
					when "00100010110" => rgb <= "111110";
					when "00100010111" => rgb <= "111110";
					when "00100011000" => rgb <= "110110";
					when "00100011001" => rgb <= "110110";
					when "00100100000" => rgb <= "101010";
					when "00100100001" => rgb <= "101010";
					when "00100100010" => rgb <= "101010";
					when "00100100011" => rgb <= "101010";
					when "00100100100" => rgb <= "101010";
					when "00100100101" => rgb <= "101010";
					when "00100100110" => rgb <= "111110";
					when "00100100111" => rgb <= "111110";
					when "00100101000" => rgb <= "111110";
					when "00100101001" => rgb <= "111110";
					when "00100101010" => rgb <= "111110";
					when "00100101011" => rgb <= "111110";
					when "00100101100" => rgb <= "111110";
					when "00100101101" => rgb <= "111110";
					when "00100101110" => rgb <= "111110";
					when "00100101111" => rgb <= "111110";
					when "00100110000" => rgb <= "111110";
					when "00100110001" => rgb <= "111110";
					when "00100110010" => rgb <= "111110";
					when "00100110011" => rgb <= "111110";
					when "00100110100" => rgb <= "111110";
					when "00100110101" => rgb <= "111110";
					when "00100110110" => rgb <= "111110";
					when "00100110111" => rgb <= "111110";
					when "00100111000" => rgb <= "110110";
					when "00100111001" => rgb <= "110110";
					when "00101000000" => rgb <= "101010";
					when "00101000001" => rgb <= "101010";
					when "00101000010" => rgb <= "101010";
					when "00101000011" => rgb <= "101010";
					when "00101000100" => rgb <= "111110";
					when "00101000101" => rgb <= "111110";
					when "00101000110" => rgb <= "111110";
					when "00101000111" => rgb <= "111110";
					when "00101001000" => rgb <= "111110";
					when "00101001001" => rgb <= "111110";
					when "00101001010" => rgb <= "111110";
					when "00101001011" => rgb <= "111110";
					when "00101001100" => rgb <= "111110";
					when "00101001101" => rgb <= "111110";
					when "00101001110" => rgb <= "111110";
					when "00101001111" => rgb <= "111110";
					when "00101010000" => rgb <= "111110";
					when "00101010001" => rgb <= "111110";
					when "00101010010" => rgb <= "111110";
					when "00101010011" => rgb <= "111110";
					when "00101010100" => rgb <= "111110";
					when "00101010101" => rgb <= "111110";
					when "00101010110" => rgb <= "111110";
					when "00101010111" => rgb <= "111110";
					when "00101011000" => rgb <= "110110";
					when "00101011001" => rgb <= "110110";
					when "00101100000" => rgb <= "101010";
					when "00101100001" => rgb <= "101010";
					when "00101100010" => rgb <= "101010";
					when "00101100011" => rgb <= "101010";
					when "00101100100" => rgb <= "111110";
					when "00101100101" => rgb <= "111110";
					when "00101100110" => rgb <= "111110";
					when "00101100111" => rgb <= "111110";
					when "00101101000" => rgb <= "111110";
					when "00101101001" => rgb <= "111110";
					when "00101101010" => rgb <= "111110";
					when "00101101011" => rgb <= "111110";
					when "00101101100" => rgb <= "111110";
					when "00101101101" => rgb <= "111110";
					when "00101101110" => rgb <= "111110";
					when "00101101111" => rgb <= "111110";
					when "00101110000" => rgb <= "111110";
					when "00101110001" => rgb <= "111110";
					when "00101110010" => rgb <= "111110";
					when "00101110011" => rgb <= "111110";
					when "00101110100" => rgb <= "111110";
					when "00101110101" => rgb <= "111110";
					when "00101110110" => rgb <= "111110";
					when "00101110111" => rgb <= "111110";
					when "00101111000" => rgb <= "110110";
					when "00101111001" => rgb <= "110110";
					when "00110000000" => rgb <= "101010";
					when "00110000001" => rgb <= "101010";
					when "00110000010" => rgb <= "101010";
					when "00110000011" => rgb <= "101010";
					when "00110000100" => rgb <= "111110";
					when "00110000101" => rgb <= "111110";
					when "00110000110" => rgb <= "111110";
					when "00110000111" => rgb <= "111110";
					when "00110001000" => rgb <= "000000";
					when "00110001001" => rgb <= "000000";
					when "00110001010" => rgb <= "111110";
					when "00110001011" => rgb <= "111110";
					when "00110001100" => rgb <= "111110";
					when "00110001101" => rgb <= "111110";
					when "00110001110" => rgb <= "111110";
					when "00110001111" => rgb <= "111110";
					when "00110010000" => rgb <= "111110";
					when "00110010001" => rgb <= "111110";
					when "00110010010" => rgb <= "111110";
					when "00110010011" => rgb <= "111110";
					when "00110010100" => rgb <= "111110";
					when "00110010101" => rgb <= "111110";
					when "00110010110" => rgb <= "111110";
					when "00110010111" => rgb <= "111110";
					when "00110011000" => rgb <= "110110";
					when "00110011001" => rgb <= "110110";
					when "00110100000" => rgb <= "101010";
					when "00110100001" => rgb <= "101010";
					when "00110100010" => rgb <= "101010";
					when "00110100011" => rgb <= "101010";
					when "00110100100" => rgb <= "111110";
					when "00110100101" => rgb <= "111110";
					when "00110100110" => rgb <= "111110";
					when "00110100111" => rgb <= "111110";
					when "00110101000" => rgb <= "000000";
					when "00110101001" => rgb <= "000000";
					when "00110101010" => rgb <= "111110";
					when "00110101011" => rgb <= "111110";
					when "00110101100" => rgb <= "111110";
					when "00110101101" => rgb <= "111110";
					when "00110101110" => rgb <= "111110";
					when "00110101111" => rgb <= "111110";
					when "00110110000" => rgb <= "111110";
					when "00110110001" => rgb <= "111110";
					when "00110110010" => rgb <= "111110";
					when "00110110011" => rgb <= "111110";
					when "00110110100" => rgb <= "111110";
					when "00110110101" => rgb <= "111110";
					when "00110110110" => rgb <= "111110";
					when "00110110111" => rgb <= "111110";
					when "00110111000" => rgb <= "110110";
					when "00110111001" => rgb <= "110110";
					when "00111000000" => rgb <= "101010";
					when "00111000001" => rgb <= "101010";
					when "00111000010" => rgb <= "101010";
					when "00111000011" => rgb <= "101010";
					when "00111000100" => rgb <= "111110";
					when "00111000101" => rgb <= "111110";
					when "00111000110" => rgb <= "000000";
					when "00111000111" => rgb <= "000000";
					when "00111001000" => rgb <= "111001";
					when "00111001001" => rgb <= "111001";
					when "00111001010" => rgb <= "000000";
					when "00111001011" => rgb <= "000000";
					when "00111001100" => rgb <= "111110";
					when "00111001101" => rgb <= "111110";
					when "00111001110" => rgb <= "111110";
					when "00111001111" => rgb <= "111110";
					when "00111010000" => rgb <= "111110";
					when "00111010001" => rgb <= "111110";
					when "00111010010" => rgb <= "000000";
					when "00111010011" => rgb <= "000000";
					when "00111010100" => rgb <= "000000";
					when "00111010101" => rgb <= "000000";
					when "00111010110" => rgb <= "111110";
					when "00111010111" => rgb <= "111110";
					when "00111011000" => rgb <= "110110";
					when "00111011001" => rgb <= "110110";
					when "00111100000" => rgb <= "101010";
					when "00111100001" => rgb <= "101010";
					when "00111100010" => rgb <= "101010";
					when "00111100011" => rgb <= "101010";
					when "00111100100" => rgb <= "111110";
					when "00111100101" => rgb <= "111110";
					when "00111100110" => rgb <= "000000";
					when "00111100111" => rgb <= "000000";
					when "00111101000" => rgb <= "111001";
					when "00111101001" => rgb <= "111001";
					when "00111101010" => rgb <= "000000";
					when "00111101011" => rgb <= "000000";
					when "00111101100" => rgb <= "111110";
					when "00111101101" => rgb <= "111110";
					when "00111101110" => rgb <= "111110";
					when "00111101111" => rgb <= "111110";
					when "00111110000" => rgb <= "111110";
					when "00111110001" => rgb <= "111110";
					when "00111110010" => rgb <= "000000";
					when "00111110011" => rgb <= "000000";
					when "00111110100" => rgb <= "000000";
					when "00111110101" => rgb <= "000000";
					when "00111110110" => rgb <= "111110";
					when "00111110111" => rgb <= "111110";
					when "00111111000" => rgb <= "110110";
					when "00111111001" => rgb <= "110110";
					when "01000000000" => rgb <= "101010";
					when "01000000001" => rgb <= "101010";
					when "01000000010" => rgb <= "101010";
					when "01000000011" => rgb <= "101010";
					when "01000000100" => rgb <= "111110";
					when "01000000101" => rgb <= "111110";
					when "01000000110" => rgb <= "111001";
					when "01000000111" => rgb <= "111001";
					when "01000001000" => rgb <= "111110";
					when "01000001001" => rgb <= "111110";
					when "01000001010" => rgb <= "111001";
					when "01000001011" => rgb <= "111001";
					when "01000001100" => rgb <= "000000";
					when "01000001101" => rgb <= "000000";
					when "01000001110" => rgb <= "000000";
					when "01000001111" => rgb <= "000000";
					when "01000010000" => rgb <= "000000";
					when "01000010001" => rgb <= "000000";
					when "01000010010" => rgb <= "111110";
					when "01000010011" => rgb <= "111110";
					when "01000010100" => rgb <= "101010";
					when "01000010101" => rgb <= "101010";
					when "01000010110" => rgb <= "000000";
					when "01000010111" => rgb <= "000000";
					when "01000011000" => rgb <= "110110";
					when "01000011001" => rgb <= "110110";
					when "01000100000" => rgb <= "101010";
					when "01000100001" => rgb <= "101010";
					when "01000100010" => rgb <= "101010";
					when "01000100011" => rgb <= "101010";
					when "01000100100" => rgb <= "111110";
					when "01000100101" => rgb <= "111110";
					when "01000100110" => rgb <= "111001";
					when "01000100111" => rgb <= "111001";
					when "01000101000" => rgb <= "111110";
					when "01000101001" => rgb <= "111110";
					when "01000101010" => rgb <= "111001";
					when "01000101011" => rgb <= "111001";
					when "01000101100" => rgb <= "000000";
					when "01000101101" => rgb <= "000000";
					when "01000101110" => rgb <= "000000";
					when "01000101111" => rgb <= "000000";
					when "01000110000" => rgb <= "000000";
					when "01000110001" => rgb <= "000000";
					when "01000110010" => rgb <= "111110";
					when "01000110011" => rgb <= "111110";
					when "01000110100" => rgb <= "101010";
					when "01000110101" => rgb <= "101010";
					when "01000110110" => rgb <= "000000";
					when "01000110111" => rgb <= "000000";
					when "01000111000" => rgb <= "110110";
					when "01000111001" => rgb <= "110110";
					when "01001000000" => rgb <= "101010";
					when "01001000001" => rgb <= "101010";
					when "01001000010" => rgb <= "101010";
					when "01001000011" => rgb <= "101010";
					when "01001000100" => rgb <= "111110";
					when "01001000101" => rgb <= "111110";
					when "01001000110" => rgb <= "111001";
					when "01001000111" => rgb <= "111001";
					when "01001001000" => rgb <= "111110";
					when "01001001001" => rgb <= "111110";
					when "01001001010" => rgb <= "111110";
					when "01001001011" => rgb <= "111110";
					when "01001001100" => rgb <= "111110";
					when "01001001101" => rgb <= "111110";
					when "01001001110" => rgb <= "111110";
					when "01001001111" => rgb <= "111110";
					when "01001010000" => rgb <= "111110";
					when "01001010001" => rgb <= "111110";
					when "01001010010" => rgb <= "000000";
					when "01001010011" => rgb <= "000000";
					when "01001010100" => rgb <= "000000";
					when "01001010101" => rgb <= "000000";
					when "01001010110" => rgb <= "111110";
					when "01001010111" => rgb <= "111110";
					when "01001011000" => rgb <= "111001";
					when "01001011001" => rgb <= "111001";
					when "01001100000" => rgb <= "101010";
					when "01001100001" => rgb <= "101010";
					when "01001100010" => rgb <= "101010";
					when "01001100011" => rgb <= "101010";
					when "01001100100" => rgb <= "111110";
					when "01001100101" => rgb <= "111110";
					when "01001100110" => rgb <= "111001";
					when "01001100111" => rgb <= "111001";
					when "01001101000" => rgb <= "111110";
					when "01001101001" => rgb <= "111110";
					when "01001101010" => rgb <= "111110";
					when "01001101011" => rgb <= "111110";
					when "01001101100" => rgb <= "111110";
					when "01001101101" => rgb <= "111110";
					when "01001101110" => rgb <= "111110";
					when "01001101111" => rgb <= "111110";
					when "01001110000" => rgb <= "111110";
					when "01001110001" => rgb <= "111110";
					when "01001110010" => rgb <= "000000";
					when "01001110011" => rgb <= "000000";
					when "01001110100" => rgb <= "000000";
					when "01001110101" => rgb <= "000000";
					when "01001110110" => rgb <= "111110";
					when "01001110111" => rgb <= "111110";
					when "01001111000" => rgb <= "111001";
					when "01001111001" => rgb <= "111001";
					when "01010000000" => rgb <= "101010";
					when "01010000001" => rgb <= "101010";
					when "01010000010" => rgb <= "101010";
					when "01010000011" => rgb <= "101010";
					when "01010000100" => rgb <= "111110";
					when "01010000101" => rgb <= "111110";
					when "01010000110" => rgb <= "111001";
					when "01010000111" => rgb <= "111001";
					when "01010001000" => rgb <= "111110";
					when "01010001001" => rgb <= "111110";
					when "01010001010" => rgb <= "111110";
					when "01010001011" => rgb <= "111110";
					when "01010001100" => rgb <= "111110";
					when "01010001101" => rgb <= "111110";
					when "01010001110" => rgb <= "111110";
					when "01010001111" => rgb <= "111110";
					when "01010010000" => rgb <= "111110";
					when "01010010001" => rgb <= "111110";
					when "01010010010" => rgb <= "111110";
					when "01010010011" => rgb <= "111110";
					when "01010010100" => rgb <= "111001";
					when "01010010101" => rgb <= "111001";
					when "01010010110" => rgb <= "111110";
					when "01010010111" => rgb <= "111110";
					when "01010011000" => rgb <= "111001";
					when "01010011001" => rgb <= "111001";
					when "01010100000" => rgb <= "101010";
					when "01010100001" => rgb <= "101010";
					when "01010100010" => rgb <= "101010";
					when "01010100011" => rgb <= "101010";
					when "01010100100" => rgb <= "111110";
					when "01010100101" => rgb <= "111110";
					when "01010100110" => rgb <= "111001";
					when "01010100111" => rgb <= "111001";
					when "01010101000" => rgb <= "111110";
					when "01010101001" => rgb <= "111110";
					when "01010101010" => rgb <= "111110";
					when "01010101011" => rgb <= "111110";
					when "01010101100" => rgb <= "111110";
					when "01010101101" => rgb <= "111110";
					when "01010101110" => rgb <= "111110";
					when "01010101111" => rgb <= "111110";
					when "01010110000" => rgb <= "111110";
					when "01010110001" => rgb <= "111110";
					when "01010110010" => rgb <= "111110";
					when "01010110011" => rgb <= "111110";
					when "01010110100" => rgb <= "111001";
					when "01010110101" => rgb <= "111001";
					when "01010110110" => rgb <= "111110";
					when "01010110111" => rgb <= "111110";
					when "01010111000" => rgb <= "111001";
					when "01010111001" => rgb <= "111001";
					when "01011000000" => rgb <= "101010";
					when "01011000001" => rgb <= "101010";
					when "01011000010" => rgb <= "101010";
					when "01011000011" => rgb <= "101010";
					when "01011000100" => rgb <= "111110";
					when "01011000101" => rgb <= "111110";
					when "01011000110" => rgb <= "111001";
					when "01011000111" => rgb <= "111001";
					when "01011001000" => rgb <= "111110";
					when "01011001001" => rgb <= "111110";
					when "01011001010" => rgb <= "111001";
					when "01011001011" => rgb <= "111001";
					when "01011001100" => rgb <= "111110";
					when "01011001101" => rgb <= "111110";
					when "01011001110" => rgb <= "111110";
					when "01011001111" => rgb <= "111110";
					when "01011010000" => rgb <= "111110";
					when "01011010001" => rgb <= "111110";
					when "01011010010" => rgb <= "111110";
					when "01011010011" => rgb <= "111110";
					when "01011010100" => rgb <= "111001";
					when "01011010101" => rgb <= "111001";
					when "01011010110" => rgb <= "111110";
					when "01011010111" => rgb <= "111110";
					when "01011011000" => rgb <= "111001";
					when "01011011001" => rgb <= "111001";
					when "01011100000" => rgb <= "101010";
					when "01011100001" => rgb <= "101010";
					when "01011100010" => rgb <= "101010";
					when "01011100011" => rgb <= "101010";
					when "01011100100" => rgb <= "111110";
					when "01011100101" => rgb <= "111110";
					when "01011100110" => rgb <= "111001";
					when "01011100111" => rgb <= "111001";
					when "01011101000" => rgb <= "111110";
					when "01011101001" => rgb <= "111110";
					when "01011101010" => rgb <= "111001";
					when "01011101011" => rgb <= "111001";
					when "01011101100" => rgb <= "111110";
					when "01011101101" => rgb <= "111110";
					when "01011101110" => rgb <= "111110";
					when "01011101111" => rgb <= "111110";
					when "01011110000" => rgb <= "111110";
					when "01011110001" => rgb <= "111110";
					when "01011110010" => rgb <= "111110";
					when "01011110011" => rgb <= "111110";
					when "01011110100" => rgb <= "111001";
					when "01011110101" => rgb <= "111001";
					when "01011110110" => rgb <= "111110";
					when "01011110111" => rgb <= "111110";
					when "01011111000" => rgb <= "111001";
					when "01011111001" => rgb <= "111001";
					when "01100000000" => rgb <= "101010";
					when "01100000001" => rgb <= "101010";
					when "01100000010" => rgb <= "101010";
					when "01100000011" => rgb <= "101010";
					when "01100000100" => rgb <= "111110";
					when "01100000101" => rgb <= "111110";
					when "01100000110" => rgb <= "111110";
					when "01100000111" => rgb <= "111110";
					when "01100001000" => rgb <= "111001";
					when "01100001001" => rgb <= "111001";
					when "01100001010" => rgb <= "111110";
					when "01100001011" => rgb <= "111110";
					when "01100001100" => rgb <= "111110";
					when "01100001101" => rgb <= "111110";
					when "01100001110" => rgb <= "111110";
					when "01100001111" => rgb <= "111110";
					when "01100010000" => rgb <= "111110";
					when "01100010001" => rgb <= "111110";
					when "01100010010" => rgb <= "111001";
					when "01100010011" => rgb <= "111001";
					when "01100010100" => rgb <= "111110";
					when "01100010101" => rgb <= "111110";
					when "01100010110" => rgb <= "111110";
					when "01100010111" => rgb <= "111110";
					when "01100011000" => rgb <= "111001";
					when "01100011001" => rgb <= "111001";
					when "01100100000" => rgb <= "101010";
					when "01100100001" => rgb <= "101010";
					when "01100100010" => rgb <= "101010";
					when "01100100011" => rgb <= "101010";
					when "01100100100" => rgb <= "111110";
					when "01100100101" => rgb <= "111110";
					when "01100100110" => rgb <= "111110";
					when "01100100111" => rgb <= "111110";
					when "01100101000" => rgb <= "111001";
					when "01100101001" => rgb <= "111001";
					when "01100101010" => rgb <= "111110";
					when "01100101011" => rgb <= "111110";
					when "01100101100" => rgb <= "111110";
					when "01100101101" => rgb <= "111110";
					when "01100101110" => rgb <= "111110";
					when "01100101111" => rgb <= "111110";
					when "01100110000" => rgb <= "111110";
					when "01100110001" => rgb <= "111110";
					when "01100110010" => rgb <= "111001";
					when "01100110011" => rgb <= "111001";
					when "01100110100" => rgb <= "111110";
					when "01100110101" => rgb <= "111110";
					when "01100110110" => rgb <= "111110";
					when "01100110111" => rgb <= "111110";
					when "01100111000" => rgb <= "111001";
					when "01100111001" => rgb <= "111001";
					when "01101000000" => rgb <= "101010";
					when "01101000001" => rgb <= "101010";
					when "01101000010" => rgb <= "101010";
					when "01101000011" => rgb <= "101010";
					when "01101000100" => rgb <= "111110";
					when "01101000101" => rgb <= "111110";
					when "01101000110" => rgb <= "111110";
					when "01101000111" => rgb <= "111110";
					when "01101001000" => rgb <= "111110";
					when "01101001001" => rgb <= "111110";
					when "01101001010" => rgb <= "111110";
					when "01101001011" => rgb <= "111110";
					when "01101001100" => rgb <= "111110";
					when "01101001101" => rgb <= "111110";
					when "01101001110" => rgb <= "111110";
					when "01101001111" => rgb <= "111110";
					when "01101010000" => rgb <= "111110";
					when "01101010001" => rgb <= "111110";
					when "01101010010" => rgb <= "111110";
					when "01101010011" => rgb <= "111110";
					when "01101010100" => rgb <= "111001";
					when "01101010101" => rgb <= "111001";
					when "01101010110" => rgb <= "111001";
					when "01101010111" => rgb <= "111001";
					when "01101011000" => rgb <= "110110";
					when "01101011001" => rgb <= "110110";
					when "01101100000" => rgb <= "101010";
					when "01101100001" => rgb <= "101010";
					when "01101100010" => rgb <= "101010";
					when "01101100011" => rgb <= "101010";
					when "01101100100" => rgb <= "111110";
					when "01101100101" => rgb <= "111110";
					when "01101100110" => rgb <= "111110";
					when "01101100111" => rgb <= "111110";
					when "01101101000" => rgb <= "111110";
					when "01101101001" => rgb <= "111110";
					when "01101101010" => rgb <= "111110";
					when "01101101011" => rgb <= "111110";
					when "01101101100" => rgb <= "111110";
					when "01101101101" => rgb <= "111110";
					when "01101101110" => rgb <= "111110";
					when "01101101111" => rgb <= "111110";
					when "01101110000" => rgb <= "111110";
					when "01101110001" => rgb <= "111110";
					when "01101110010" => rgb <= "111110";
					when "01101110011" => rgb <= "111110";
					when "01101110100" => rgb <= "111001";
					when "01101110101" => rgb <= "111001";
					when "01101110110" => rgb <= "111001";
					when "01101110111" => rgb <= "111001";
					when "01101111000" => rgb <= "110110";
					when "01101111001" => rgb <= "110110";
					when "01110000000" => rgb <= "101010";
					when "01110000001" => rgb <= "101010";
					when "01110000010" => rgb <= "101010";
					when "01110000011" => rgb <= "101010";
					when "01110000100" => rgb <= "111110";
					when "01110000101" => rgb <= "111110";
					when "01110000110" => rgb <= "111110";
					when "01110000111" => rgb <= "111110";
					when "01110001000" => rgb <= "111110";
					when "01110001001" => rgb <= "111110";
					when "01110001010" => rgb <= "111110";
					when "01110001011" => rgb <= "111110";
					when "01110001100" => rgb <= "111110";
					when "01110001101" => rgb <= "111110";
					when "01110001110" => rgb <= "111110";
					when "01110001111" => rgb <= "111110";
					when "01110010000" => rgb <= "111110";
					when "01110010001" => rgb <= "111110";
					when "01110010010" => rgb <= "111110";
					when "01110010011" => rgb <= "111110";
					when "01110010100" => rgb <= "111110";
					when "01110010101" => rgb <= "111110";
					when "01110010110" => rgb <= "111110";
					when "01110010111" => rgb <= "111110";
					when "01110011000" => rgb <= "110110";
					when "01110011001" => rgb <= "110110";
					when "01110100000" => rgb <= "101010";
					when "01110100001" => rgb <= "101010";
					when "01110100010" => rgb <= "101010";
					when "01110100011" => rgb <= "101010";
					when "01110100100" => rgb <= "111110";
					when "01110100101" => rgb <= "111110";
					when "01110100110" => rgb <= "111110";
					when "01110100111" => rgb <= "111110";
					when "01110101000" => rgb <= "111110";
					when "01110101001" => rgb <= "111110";
					when "01110101010" => rgb <= "111110";
					when "01110101011" => rgb <= "111110";
					when "01110101100" => rgb <= "111110";
					when "01110101101" => rgb <= "111110";
					when "01110101110" => rgb <= "111110";
					when "01110101111" => rgb <= "111110";
					when "01110110000" => rgb <= "111110";
					when "01110110001" => rgb <= "111110";
					when "01110110010" => rgb <= "111110";
					when "01110110011" => rgb <= "111110";
					when "01110110100" => rgb <= "111110";
					when "01110110101" => rgb <= "111110";
					when "01110110110" => rgb <= "111110";
					when "01110110111" => rgb <= "111110";
					when "01110111000" => rgb <= "110110";
					when "01110111001" => rgb <= "110110";
					when "01111000000" => rgb <= "101010";
					when "01111000001" => rgb <= "101010";
					when "01111000010" => rgb <= "111110";
					when "01111000011" => rgb <= "111110";
					when "01111000100" => rgb <= "111110";
					when "01111000101" => rgb <= "111110";
					when "01111000110" => rgb <= "111110";
					when "01111000111" => rgb <= "111110";
					when "01111001000" => rgb <= "111110";
					when "01111001001" => rgb <= "111110";
					when "01111001010" => rgb <= "111110";
					when "01111001011" => rgb <= "111110";
					when "01111001100" => rgb <= "111110";
					when "01111001101" => rgb <= "111110";
					when "01111001110" => rgb <= "111110";
					when "01111001111" => rgb <= "111110";
					when "01111010000" => rgb <= "110101";
					when "01111010001" => rgb <= "110101";
					when "01111010010" => rgb <= "110101";
					when "01111010011" => rgb <= "110101";
					when "01111010100" => rgb <= "110101";
					when "01111010101" => rgb <= "110101";
					when "01111010110" => rgb <= "110101";
					when "01111010111" => rgb <= "110101";
					when "01111011000" => rgb <= "110110";
					when "01111011001" => rgb <= "110110";
					when "01111100000" => rgb <= "101010";
					when "01111100001" => rgb <= "101010";
					when "01111100010" => rgb <= "111110";
					when "01111100011" => rgb <= "111110";
					when "01111100100" => rgb <= "111110";
					when "01111100101" => rgb <= "111110";
					when "01111100110" => rgb <= "111110";
					when "01111100111" => rgb <= "111110";
					when "01111101000" => rgb <= "111110";
					when "01111101001" => rgb <= "111110";
					when "01111101010" => rgb <= "111110";
					when "01111101011" => rgb <= "111110";
					when "01111101100" => rgb <= "111110";
					when "01111101101" => rgb <= "111110";
					when "01111101110" => rgb <= "111110";
					when "01111101111" => rgb <= "111110";
					when "01111110000" => rgb <= "110101";
					when "01111110001" => rgb <= "110101";
					when "01111110010" => rgb <= "110101";
					when "01111110011" => rgb <= "110101";
					when "01111110100" => rgb <= "110101";
					when "01111110101" => rgb <= "110101";
					when "01111110110" => rgb <= "110101";
					when "01111110111" => rgb <= "110101";
					when "01111111000" => rgb <= "110110";
					when "01111111001" => rgb <= "110110";
					when "10000000000" => rgb <= "101010";
					when "10000000001" => rgb <= "101010";
					when "10000000010" => rgb <= "111110";
					when "10000000011" => rgb <= "111110";
					when "10000000100" => rgb <= "111110";
					when "10000000101" => rgb <= "111110";
					when "10000000110" => rgb <= "111110";
					when "10000000111" => rgb <= "111110";
					when "10000001000" => rgb <= "111110";
					when "10000001001" => rgb <= "111110";
					when "10000001010" => rgb <= "111110";
					when "10000001011" => rgb <= "111110";
					when "10000001100" => rgb <= "111110";
					when "10000001101" => rgb <= "111110";
					when "10000001110" => rgb <= "111110";
					when "10000001111" => rgb <= "111110";
					when "10000010000" => rgb <= "110101";
					when "10000010001" => rgb <= "110101";
					when "10000010010" => rgb <= "111111";
					when "10000010011" => rgb <= "111111";
					when "10000010100" => rgb <= "111111";
					when "10000010101" => rgb <= "111111";
					when "10000010110" => rgb <= "111111";
					when "10000010111" => rgb <= "111111";
					when "10000011000" => rgb <= "110110";
					when "10000011001" => rgb <= "110110";
					when "10000100000" => rgb <= "101010";
					when "10000100001" => rgb <= "101010";
					when "10000100010" => rgb <= "111110";
					when "10000100011" => rgb <= "111110";
					when "10000100100" => rgb <= "111110";
					when "10000100101" => rgb <= "111110";
					when "10000100110" => rgb <= "111110";
					when "10000100111" => rgb <= "111110";
					when "10000101000" => rgb <= "111110";
					when "10000101001" => rgb <= "111110";
					when "10000101010" => rgb <= "111110";
					when "10000101011" => rgb <= "111110";
					when "10000101100" => rgb <= "111110";
					when "10000101101" => rgb <= "111110";
					when "10000101110" => rgb <= "111110";
					when "10000101111" => rgb <= "111110";
					when "10000110000" => rgb <= "110101";
					when "10000110001" => rgb <= "110101";
					when "10000110010" => rgb <= "111111";
					when "10000110011" => rgb <= "111111";
					when "10000110100" => rgb <= "111111";
					when "10000110101" => rgb <= "111111";
					when "10000110110" => rgb <= "111111";
					when "10000110111" => rgb <= "111111";
					when "10000111000" => rgb <= "110110";
					when "10000111001" => rgb <= "110110";
					when "10001000000" => rgb <= "110110";
					when "10001000001" => rgb <= "110110";
					when "10001000010" => rgb <= "111110";
					when "10001000011" => rgb <= "111110";
					when "10001000100" => rgb <= "111110";
					when "10001000101" => rgb <= "111110";
					when "10001000110" => rgb <= "111110";
					when "10001000111" => rgb <= "111110";
					when "10001001000" => rgb <= "111110";
					when "10001001001" => rgb <= "111110";
					when "10001001010" => rgb <= "111110";
					when "10001001011" => rgb <= "111110";
					when "10001001100" => rgb <= "111110";
					when "10001001101" => rgb <= "111110";
					when "10001001110" => rgb <= "111110";
					when "10001001111" => rgb <= "111110";
					when "10001010000" => rgb <= "111110";
					when "10001010001" => rgb <= "111110";
					when "10001010010" => rgb <= "110101";
					when "10001010011" => rgb <= "110101";
					when "10001010100" => rgb <= "110101";
					when "10001010101" => rgb <= "110101";
					when "10001010110" => rgb <= "110101";
					when "10001010111" => rgb <= "110101";
					when "10001011000" => rgb <= "110110";
					when "10001011001" => rgb <= "110110";
					when "10001100000" => rgb <= "110110";
					when "10001100001" => rgb <= "110110";
					when "10001100010" => rgb <= "111110";
					when "10001100011" => rgb <= "111110";
					when "10001100100" => rgb <= "111110";
					when "10001100101" => rgb <= "111110";
					when "10001100110" => rgb <= "111110";
					when "10001100111" => rgb <= "111110";
					when "10001101000" => rgb <= "111110";
					when "10001101001" => rgb <= "111110";
					when "10001101010" => rgb <= "111110";
					when "10001101011" => rgb <= "111110";
					when "10001101100" => rgb <= "111110";
					when "10001101101" => rgb <= "111110";
					when "10001101110" => rgb <= "111110";
					when "10001101111" => rgb <= "111110";
					when "10001110000" => rgb <= "111110";
					when "10001110001" => rgb <= "111110";
					when "10001110010" => rgb <= "110101";
					when "10001110011" => rgb <= "110101";
					when "10001110100" => rgb <= "110101";
					when "10001110101" => rgb <= "110101";
					when "10001110110" => rgb <= "110101";
					when "10001110111" => rgb <= "110101";
					when "10001111000" => rgb <= "110110";
					when "10001111001" => rgb <= "110110";
					when "10010000000" => rgb <= "110110";
					when "10010000001" => rgb <= "110110";
					when "10010000010" => rgb <= "110110";
					when "10010000011" => rgb <= "110110";
					when "10010000100" => rgb <= "111110";
					when "10010000101" => rgb <= "111110";
					when "10010000110" => rgb <= "111110";
					when "10010000111" => rgb <= "111110";
					when "10010001000" => rgb <= "111110";
					when "10010001001" => rgb <= "111110";
					when "10010001010" => rgb <= "111110";
					when "10010001011" => rgb <= "111110";
					when "10010001100" => rgb <= "111110";
					when "10010001101" => rgb <= "111110";
					when "10010001110" => rgb <= "111110";
					when "10010001111" => rgb <= "111110";
					when "10010010000" => rgb <= "111110";
					when "10010010001" => rgb <= "111110";
					when "10010010010" => rgb <= "111110";
					when "10010010011" => rgb <= "111110";
					when "10010010100" => rgb <= "111110";
					when "10010010101" => rgb <= "111110";
					when "10010010110" => rgb <= "111110";
					when "10010010111" => rgb <= "111110";
					when "10010011000" => rgb <= "110110";
					when "10010011001" => rgb <= "110110";
					when "10010100000" => rgb <= "110110";
					when "10010100001" => rgb <= "110110";
					when "10010100010" => rgb <= "110110";
					when "10010100011" => rgb <= "110110";
					when "10010100100" => rgb <= "111110";
					when "10010100101" => rgb <= "111110";
					when "10010100110" => rgb <= "111110";
					when "10010100111" => rgb <= "111110";
					when "10010101000" => rgb <= "111110";
					when "10010101001" => rgb <= "111110";
					when "10010101010" => rgb <= "111110";
					when "10010101011" => rgb <= "111110";
					when "10010101100" => rgb <= "111110";
					when "10010101101" => rgb <= "111110";
					when "10010101110" => rgb <= "111110";
					when "10010101111" => rgb <= "111110";
					when "10010110000" => rgb <= "111110";
					when "10010110001" => rgb <= "111110";
					when "10010110010" => rgb <= "111110";
					when "10010110011" => rgb <= "111110";
					when "10010110100" => rgb <= "111110";
					when "10010110101" => rgb <= "111110";
					when "10010110110" => rgb <= "111110";
					when "10010110111" => rgb <= "111110";
					when "10010111000" => rgb <= "110110";
					when "10010111001" => rgb <= "110110";
					when "10011000000" => rgb <= "110110";
					when "10011000001" => rgb <= "110110";
					when "10011000010" => rgb <= "110110";
					when "10011000011" => rgb <= "110110";
					when "10011000100" => rgb <= "000110";
					when "10011000101" => rgb <= "000110";
					when "10011000110" => rgb <= "000110";
					when "10011000111" => rgb <= "000110";
					when "10011001000" => rgb <= "000110";
					when "10011001001" => rgb <= "000110";
					when "10011001010" => rgb <= "000110";
					when "10011001011" => rgb <= "000110";
					when "10011001100" => rgb <= "000110";
					when "10011001101" => rgb <= "000110";
					when "10011001110" => rgb <= "000110";
					when "10011001111" => rgb <= "000110";
					when "10011010000" => rgb <= "000110";
					when "10011010001" => rgb <= "000110";
					when "10011010010" => rgb <= "111111";
					when "10011010011" => rgb <= "111111";
					when "10011010100" => rgb <= "111110";
					when "10011010101" => rgb <= "111110";
					when "10011010110" => rgb <= "111110";
					when "10011010111" => rgb <= "111110";
					when "10011011000" => rgb <= "110110";
					when "10011011001" => rgb <= "110110";
					when "10011100000" => rgb <= "110110";
					when "10011100001" => rgb <= "110110";
					when "10011100010" => rgb <= "110110";
					when "10011100011" => rgb <= "110110";
					when "10011100100" => rgb <= "000110";
					when "10011100101" => rgb <= "000110";
					when "10011100110" => rgb <= "000110";
					when "10011100111" => rgb <= "000110";
					when "10011101000" => rgb <= "000110";
					when "10011101001" => rgb <= "000110";
					when "10011101010" => rgb <= "000110";
					when "10011101011" => rgb <= "000110";
					when "10011101100" => rgb <= "000110";
					when "10011101101" => rgb <= "000110";
					when "10011101110" => rgb <= "000110";
					when "10011101111" => rgb <= "000110";
					when "10011110000" => rgb <= "000110";
					when "10011110001" => rgb <= "000110";
					when "10011110010" => rgb <= "111111";
					when "10011110011" => rgb <= "111111";
					when "10011110100" => rgb <= "111110";
					when "10011110101" => rgb <= "111110";
					when "10011110110" => rgb <= "111110";
					when "10011110111" => rgb <= "111110";
					when "10011111000" => rgb <= "110110";
					when "10011111001" => rgb <= "110110";
					when "10100000000" => rgb <= "110110";
					when "10100000001" => rgb <= "110110";
					when "10100000010" => rgb <= "110110";
					when "10100000011" => rgb <= "110110";
					when "10100000100" => rgb <= "000110";
					when "10100000101" => rgb <= "000110";
					when "10100000110" => rgb <= "000110";
					when "10100000111" => rgb <= "000110";
					when "10100001000" => rgb <= "000110";
					when "10100001001" => rgb <= "000110";
					when "10100001010" => rgb <= "000110";
					when "10100001011" => rgb <= "000110";
					when "10100001100" => rgb <= "000110";
					when "10100001101" => rgb <= "000110";
					when "10100001110" => rgb <= "000110";
					when "10100001111" => rgb <= "000110";
					when "10100010000" => rgb <= "000110";
					when "10100010001" => rgb <= "000110";
					when "10100010010" => rgb <= "000110";
					when "10100010011" => rgb <= "000110";
					when "10100010100" => rgb <= "000110";
					when "10100010101" => rgb <= "000110";
					when "10100010110" => rgb <= "111110";
					when "10100010111" => rgb <= "111110";
					when "10100011000" => rgb <= "111110";
					when "10100011001" => rgb <= "111110";
					when "10100100000" => rgb <= "110110";
					when "10100100001" => rgb <= "110110";
					when "10100100010" => rgb <= "110110";
					when "10100100011" => rgb <= "110110";
					when "10100100100" => rgb <= "000110";
					when "10100100101" => rgb <= "000110";
					when "10100100110" => rgb <= "000110";
					when "10100100111" => rgb <= "000110";
					when "10100101000" => rgb <= "000110";
					when "10100101001" => rgb <= "000110";
					when "10100101010" => rgb <= "000110";
					when "10100101011" => rgb <= "000110";
					when "10100101100" => rgb <= "000110";
					when "10100101101" => rgb <= "000110";
					when "10100101110" => rgb <= "000110";
					when "10100101111" => rgb <= "000110";
					when "10100110000" => rgb <= "000110";
					when "10100110001" => rgb <= "000110";
					when "10100110010" => rgb <= "000110";
					when "10100110011" => rgb <= "000110";
					when "10100110100" => rgb <= "000110";
					when "10100110101" => rgb <= "000110";
					when "10100110110" => rgb <= "111110";
					when "10100110111" => rgb <= "111110";
					when "10100111000" => rgb <= "111110";
					when "10100111001" => rgb <= "111110";
					when "10101000000" => rgb <= "110110";
					when "10101000001" => rgb <= "110110";
					when "10101000010" => rgb <= "110110";
					when "10101000011" => rgb <= "110110";
					when "10101000100" => rgb <= "000110";
					when "10101000101" => rgb <= "000110";
					when "10101000110" => rgb <= "000110";
					when "10101000111" => rgb <= "000110";
					when "10101001000" => rgb <= "000110";
					when "10101001001" => rgb <= "000110";
					when "10101001010" => rgb <= "000110";
					when "10101001011" => rgb <= "000110";
					when "10101001100" => rgb <= "000110";
					when "10101001101" => rgb <= "000110";
					when "10101001110" => rgb <= "000110";
					when "10101001111" => rgb <= "000110";
					when "10101010000" => rgb <= "000110";
					when "10101010001" => rgb <= "000110";
					when "10101010010" => rgb <= "000110";
					when "10101010011" => rgb <= "000110";
					when "10101010100" => rgb <= "000110";
					when "10101010101" => rgb <= "000110";
					when "10101010110" => rgb <= "111110";
					when "10101010111" => rgb <= "111110";
					when "10101011000" => rgb <= "111110";
					when "10101011001" => rgb <= "111110";
					when "10101100000" => rgb <= "110110";
					when "10101100001" => rgb <= "110110";
					when "10101100010" => rgb <= "110110";
					when "10101100011" => rgb <= "110110";
					when "10101100100" => rgb <= "000110";
					when "10101100101" => rgb <= "000110";
					when "10101100110" => rgb <= "000110";
					when "10101100111" => rgb <= "000110";
					when "10101101000" => rgb <= "000110";
					when "10101101001" => rgb <= "000110";
					when "10101101010" => rgb <= "000110";
					when "10101101011" => rgb <= "000110";
					when "10101101100" => rgb <= "000110";
					when "10101101101" => rgb <= "000110";
					when "10101101110" => rgb <= "000110";
					when "10101101111" => rgb <= "000110";
					when "10101110000" => rgb <= "000110";
					when "10101110001" => rgb <= "000110";
					when "10101110010" => rgb <= "000110";
					when "10101110011" => rgb <= "000110";
					when "10101110100" => rgb <= "000110";
					when "10101110101" => rgb <= "000110";
					when "10101110110" => rgb <= "111110";
					when "10101110111" => rgb <= "111110";
					when "10101111000" => rgb <= "111110";
					when "10101111001" => rgb <= "111110";
					when "10110000000" => rgb <= "110110";
					when "10110000001" => rgb <= "110110";
					when "10110000010" => rgb <= "110110";
					when "10110000011" => rgb <= "110110";
					when "10110000100" => rgb <= "000110";
					when "10110000101" => rgb <= "000110";
					when "10110000110" => rgb <= "000110";
					when "10110000111" => rgb <= "000110";
					when "10110001000" => rgb <= "000110";
					when "10110001001" => rgb <= "000110";
					when "10110001010" => rgb <= "000110";
					when "10110001011" => rgb <= "000110";
					when "10110001100" => rgb <= "000110";
					when "10110001101" => rgb <= "000110";
					when "10110001110" => rgb <= "000110";
					when "10110001111" => rgb <= "000110";
					when "10110010000" => rgb <= "000110";
					when "10110010001" => rgb <= "000110";
					when "10110010010" => rgb <= "000110";
					when "10110010011" => rgb <= "000110";
					when "10110010100" => rgb <= "110000";
					when "10110010101" => rgb <= "110000";
					when "10110010110" => rgb <= "110110";
					when "10110010111" => rgb <= "110110";
					when "10110011000" => rgb <= "110110";
					when "10110011001" => rgb <= "110110";
					when "10110100000" => rgb <= "110110";
					when "10110100001" => rgb <= "110110";
					when "10110100010" => rgb <= "110110";
					when "10110100011" => rgb <= "110110";
					when "10110100100" => rgb <= "000110";
					when "10110100101" => rgb <= "000110";
					when "10110100110" => rgb <= "000110";
					when "10110100111" => rgb <= "000110";
					when "10110101000" => rgb <= "000110";
					when "10110101001" => rgb <= "000110";
					when "10110101010" => rgb <= "000110";
					when "10110101011" => rgb <= "000110";
					when "10110101100" => rgb <= "000110";
					when "10110101101" => rgb <= "000110";
					when "10110101110" => rgb <= "000110";
					when "10110101111" => rgb <= "000110";
					when "10110110000" => rgb <= "000110";
					when "10110110001" => rgb <= "000110";
					when "10110110010" => rgb <= "000110";
					when "10110110011" => rgb <= "000110";
					when "10110110100" => rgb <= "110000";
					when "10110110101" => rgb <= "110000";
					when "10110110110" => rgb <= "110110";
					when "10110110111" => rgb <= "110110";
					when "10110111000" => rgb <= "110110";
					when "10110111001" => rgb <= "110110";
					when "10111000000" => rgb <= "110110";
					when "10111000001" => rgb <= "110110";
					when "10111000010" => rgb <= "110110";
					when "10111000011" => rgb <= "110110";
					when "10111000100" => rgb <= "000110";
					when "10111000101" => rgb <= "000110";
					when "10111000110" => rgb <= "000110";
					when "10111000111" => rgb <= "000110";
					when "10111001000" => rgb <= "000110";
					when "10111001001" => rgb <= "000110";
					when "10111001010" => rgb <= "000110";
					when "10111001011" => rgb <= "000110";
					when "10111001100" => rgb <= "000110";
					when "10111001101" => rgb <= "000110";
					when "10111001110" => rgb <= "000110";
					when "10111001111" => rgb <= "000110";
					when "10111010000" => rgb <= "000110";
					when "10111010001" => rgb <= "000110";
					when "10111010010" => rgb <= "111111";
					when "10111010011" => rgb <= "111111";
					when "10111010100" => rgb <= "110000";
					when "10111010101" => rgb <= "110000";
					when "10111010110" => rgb <= "110110";
					when "10111010111" => rgb <= "110110";
					when "10111011000" => rgb <= "110110";
					when "10111011001" => rgb <= "110110";
					when "10111100000" => rgb <= "110110";
					when "10111100001" => rgb <= "110110";
					when "10111100010" => rgb <= "110110";
					when "10111100011" => rgb <= "110110";
					when "10111100100" => rgb <= "000110";
					when "10111100101" => rgb <= "000110";
					when "10111100110" => rgb <= "000110";
					when "10111100111" => rgb <= "000110";
					when "10111101000" => rgb <= "000110";
					when "10111101001" => rgb <= "000110";
					when "10111101010" => rgb <= "000110";
					when "10111101011" => rgb <= "000110";
					when "10111101100" => rgb <= "000110";
					when "10111101101" => rgb <= "000110";
					when "10111101110" => rgb <= "000110";
					when "10111101111" => rgb <= "000110";
					when "10111110000" => rgb <= "000110";
					when "10111110001" => rgb <= "000110";
					when "10111110010" => rgb <= "111111";
					when "10111110011" => rgb <= "111111";
					when "10111110100" => rgb <= "110000";
					when "10111110101" => rgb <= "110000";
					when "10111110110" => rgb <= "110110";
					when "10111110111" => rgb <= "110110";
					when "10111111000" => rgb <= "110110";
					when "10111111001" => rgb <= "110110";
					when "11000000000" => rgb <= "110110";
					when "11000000001" => rgb <= "110110";
					when "11000000010" => rgb <= "110110";
					when "11000000011" => rgb <= "110110";
					when "11000000100" => rgb <= "000110";
					when "11000000101" => rgb <= "000110";
					when "11000000110" => rgb <= "000110";
					when "11000000111" => rgb <= "000110";
					when "11000001000" => rgb <= "000110";
					when "11000001001" => rgb <= "000110";
					when "11000001010" => rgb <= "000110";
					when "11000001011" => rgb <= "000110";
					when "11000001100" => rgb <= "000110";
					when "11000001101" => rgb <= "000110";
					when "11000001110" => rgb <= "000110";
					when "11000001111" => rgb <= "000110";
					when "11000010000" => rgb <= "000110";
					when "11000010001" => rgb <= "000110";
					when "11000010010" => rgb <= "111111";
					when "11000010011" => rgb <= "111111";
					when "11000010100" => rgb <= "110000";
					when "11000010101" => rgb <= "110000";
					when "11000010110" => rgb <= "110110";
					when "11000010111" => rgb <= "110110";
					when "11000011000" => rgb <= "000000";
					when "11000011001" => rgb <= "000000";
					when "11000100000" => rgb <= "110110";
					when "11000100001" => rgb <= "110110";
					when "11000100010" => rgb <= "110110";
					when "11000100011" => rgb <= "110110";
					when "11000100100" => rgb <= "000110";
					when "11000100101" => rgb <= "000110";
					when "11000100110" => rgb <= "000110";
					when "11000100111" => rgb <= "000110";
					when "11000101000" => rgb <= "000110";
					when "11000101001" => rgb <= "000110";
					when "11000101010" => rgb <= "000110";
					when "11000101011" => rgb <= "000110";
					when "11000101100" => rgb <= "000110";
					when "11000101101" => rgb <= "000110";
					when "11000101110" => rgb <= "000110";
					when "11000101111" => rgb <= "000110";
					when "11000110000" => rgb <= "000110";
					when "11000110001" => rgb <= "000110";
					when "11000110010" => rgb <= "111111";
					when "11000110011" => rgb <= "111111";
					when "11000110100" => rgb <= "110000";
					when "11000110101" => rgb <= "110000";
					when "11000110110" => rgb <= "110110";
					when "11000110111" => rgb <= "110110";
					when "11000111000" => rgb <= "000000";
					when "11000111001" => rgb <= "000000";
					when "11001000000" => rgb <= "110110";
					when "11001000001" => rgb <= "110110";
					when "11001000010" => rgb <= "110110";
					when "11001000011" => rgb <= "110110";
					when "11001000100" => rgb <= "000110";
					when "11001000101" => rgb <= "000110";
					when "11001000110" => rgb <= "000110";
					when "11001000111" => rgb <= "000110";
					when "11001001000" => rgb <= "000110";
					when "11001001001" => rgb <= "000110";
					when "11001001010" => rgb <= "000110";
					when "11001001011" => rgb <= "000110";
					when "11001001100" => rgb <= "000110";
					when "11001001101" => rgb <= "000110";
					when "11001001110" => rgb <= "000110";
					when "11001001111" => rgb <= "000110";
					when "11001010000" => rgb <= "000110";
					when "11001010001" => rgb <= "000110";
					when "11001010010" => rgb <= "111111";
					when "11001010011" => rgb <= "111111";
					when "11001010100" => rgb <= "111111";
					when "11001010101" => rgb <= "111111";
					when "11001010110" => rgb <= "000000";
					when "11001010111" => rgb <= "000000";
					when "11001011000" => rgb <= "000000";
					when "11001011001" => rgb <= "000000";
					when "11001100000" => rgb <= "110110";
					when "11001100001" => rgb <= "110110";
					when "11001100010" => rgb <= "110110";
					when "11001100011" => rgb <= "110110";
					when "11001100100" => rgb <= "000110";
					when "11001100101" => rgb <= "000110";
					when "11001100110" => rgb <= "000110";
					when "11001100111" => rgb <= "000110";
					when "11001101000" => rgb <= "000110";
					when "11001101001" => rgb <= "000110";
					when "11001101010" => rgb <= "000110";
					when "11001101011" => rgb <= "000110";
					when "11001101100" => rgb <= "000110";
					when "11001101101" => rgb <= "000110";
					when "11001101110" => rgb <= "000110";
					when "11001101111" => rgb <= "000110";
					when "11001110000" => rgb <= "000110";
					when "11001110001" => rgb <= "000110";
					when "11001110010" => rgb <= "111111";
					when "11001110011" => rgb <= "111111";
					when "11001110100" => rgb <= "111111";
					when "11001110101" => rgb <= "111111";
					when "11001110110" => rgb <= "000000";
					when "11001110111" => rgb <= "000000";
					when "11001111000" => rgb <= "000000";
					when "11001111001" => rgb <= "000000";
					when "11010000000" => rgb <= "110110";
					when "11010000001" => rgb <= "110110";
					when "11010000010" => rgb <= "110110";
					when "11010000011" => rgb <= "110110";
					when "11010000100" => rgb <= "000110";
					when "11010000101" => rgb <= "000110";
					when "11010000110" => rgb <= "000110";
					when "11010000111" => rgb <= "000110";
					when "11010001000" => rgb <= "000110";
					when "11010001001" => rgb <= "000110";
					when "11010001010" => rgb <= "000110";
					when "11010001011" => rgb <= "000110";
					when "11010001100" => rgb <= "000110";
					when "11010001101" => rgb <= "000110";
					when "11010001110" => rgb <= "000110";
					when "11010001111" => rgb <= "000110";
					when "11010010000" => rgb <= "000110";
					when "11010010001" => rgb <= "000110";
					when "11010010010" => rgb <= "000110";
					when "11010010011" => rgb <= "000110";
					when "11010010100" => rgb <= "000110";
					when "11010010101" => rgb <= "000110";
					when "11010010110" => rgb <= "000000";
					when "11010010111" => rgb <= "000000";
					when "11010011000" => rgb <= "000000";
					when "11010011001" => rgb <= "000000";
					when "11010100000" => rgb <= "110110";
					when "11010100001" => rgb <= "110110";
					when "11010100010" => rgb <= "110110";
					when "11010100011" => rgb <= "110110";
					when "11010100100" => rgb <= "000110";
					when "11010100101" => rgb <= "000110";
					when "11010100110" => rgb <= "000110";
					when "11010100111" => rgb <= "000110";
					when "11010101000" => rgb <= "000110";
					when "11010101001" => rgb <= "000110";
					when "11010101010" => rgb <= "000110";
					when "11010101011" => rgb <= "000110";
					when "11010101100" => rgb <= "000110";
					when "11010101101" => rgb <= "000110";
					when "11010101110" => rgb <= "000110";
					when "11010101111" => rgb <= "000110";
					when "11010110000" => rgb <= "000110";
					when "11010110001" => rgb <= "000110";
					when "11010110010" => rgb <= "000110";
					when "11010110011" => rgb <= "000110";
					when "11010110100" => rgb <= "000110";
					when "11010110101" => rgb <= "000110";
					when "11010110110" => rgb <= "000000";
					when "11010110111" => rgb <= "000000";
					when "11010111000" => rgb <= "000000";
					when "11010111001" => rgb <= "000000";
					when "11011000000" => rgb <= "110110";
					when "11011000001" => rgb <= "110110";
					when "11011000010" => rgb <= "000110";
					when "11011000011" => rgb <= "000110";
					when "11011000100" => rgb <= "000110";
					when "11011000101" => rgb <= "000110";
					when "11011000110" => rgb <= "000110";
					when "11011000111" => rgb <= "000110";
					when "11011001000" => rgb <= "000110";
					when "11011001001" => rgb <= "000110";
					when "11011001010" => rgb <= "110110";
					when "11011001011" => rgb <= "110110";
					when "11011001100" => rgb <= "110110";
					when "11011001101" => rgb <= "110110";
					when "11011001110" => rgb <= "000110";
					when "11011001111" => rgb <= "000110";
					when "11011010000" => rgb <= "000110";
					when "11011010001" => rgb <= "000110";
					when "11011010010" => rgb <= "000110";
					when "11011010011" => rgb <= "000110";
					when "11011010100" => rgb <= "000110";
					when "11011010101" => rgb <= "000110";
					when "11011010110" => rgb <= "000000";
					when "11011010111" => rgb <= "000000";
					when "11011011000" => rgb <= "000000";
					when "11011011001" => rgb <= "000000";
					when "11011100000" => rgb <= "110110";
					when "11011100001" => rgb <= "110110";
					when "11011100010" => rgb <= "000110";
					when "11011100011" => rgb <= "000110";
					when "11011100100" => rgb <= "000110";
					when "11011100101" => rgb <= "000110";
					when "11011100110" => rgb <= "000110";
					when "11011100111" => rgb <= "000110";
					when "11011101000" => rgb <= "000110";
					when "11011101001" => rgb <= "000110";
					when "11011101010" => rgb <= "110110";
					when "11011101011" => rgb <= "110110";
					when "11011101100" => rgb <= "110110";
					when "11011101101" => rgb <= "110110";
					when "11011101110" => rgb <= "000110";
					when "11011101111" => rgb <= "000110";
					when "11011110000" => rgb <= "000110";
					when "11011110001" => rgb <= "000110";
					when "11011110010" => rgb <= "000110";
					when "11011110011" => rgb <= "000110";
					when "11011110100" => rgb <= "000110";
					when "11011110101" => rgb <= "000110";
					when "11011110110" => rgb <= "000000";
					when "11011110111" => rgb <= "000000";
					when "11011111000" => rgb <= "000000";
					when "11011111001" => rgb <= "000000";
					when "11100000000" => rgb <= "110110";
					when "11100000001" => rgb <= "110110";
					when "11100000010" => rgb <= "000110";
					when "11100000011" => rgb <= "000110";
					when "11100000100" => rgb <= "000110";
					when "11100000101" => rgb <= "000110";
					when "11100000110" => rgb <= "000110";
					when "11100000111" => rgb <= "000110";
					when "11100001000" => rgb <= "110110";
					when "11100001001" => rgb <= "110110";
					when "11100001010" => rgb <= "110110";
					when "11100001011" => rgb <= "110110";
					when "11100001100" => rgb <= "110110";
					when "11100001101" => rgb <= "110110";
					when "11100001110" => rgb <= "110110";
					when "11100001111" => rgb <= "110110";
					when "11100010000" => rgb <= "000110";
					when "11100010001" => rgb <= "000110";
					when "11100010010" => rgb <= "000110";
					when "11100010011" => rgb <= "000110";
					when "11100010100" => rgb <= "000110";
					when "11100010101" => rgb <= "000110";
					when "11100010110" => rgb <= "000000";
					when "11100010111" => rgb <= "000000";
					when "11100011000" => rgb <= "000000";
					when "11100011001" => rgb <= "000000";
					when "11100100000" => rgb <= "110110";
					when "11100100001" => rgb <= "110110";
					when "11100100010" => rgb <= "000110";
					when "11100100011" => rgb <= "000110";
					when "11100100100" => rgb <= "000110";
					when "11100100101" => rgb <= "000110";
					when "11100100110" => rgb <= "000110";
					when "11100100111" => rgb <= "000110";
					when "11100101000" => rgb <= "110110";
					when "11100101001" => rgb <= "110110";
					when "11100101010" => rgb <= "110110";
					when "11100101011" => rgb <= "110110";
					when "11100101100" => rgb <= "110110";
					when "11100101101" => rgb <= "110110";
					when "11100101110" => rgb <= "110110";
					when "11100101111" => rgb <= "110110";
					when "11100110000" => rgb <= "000110";
					when "11100110001" => rgb <= "000110";
					when "11100110010" => rgb <= "000110";
					when "11100110011" => rgb <= "000110";
					when "11100110100" => rgb <= "000110";
					when "11100110101" => rgb <= "000110";
					when "11100110110" => rgb <= "000000";
					when "11100110111" => rgb <= "000000";
					when "11100111000" => rgb <= "000000";
					when "11100111001" => rgb <= "000000";
					when "11101000000" => rgb <= "110110";
					when "11101000001" => rgb <= "110110";
					when "11101000010" => rgb <= "000000";
					when "11101000011" => rgb <= "000000";
					when "11101000100" => rgb <= "000000";
					when "11101000101" => rgb <= "000000";
					when "11101000110" => rgb <= "000000";
					when "11101000111" => rgb <= "000000";
					when "11101001000" => rgb <= "110110";
					when "11101001001" => rgb <= "110110";
					when "11101001010" => rgb <= "110110";
					when "11101001011" => rgb <= "110110";
					when "11101001100" => rgb <= "110110";
					when "11101001101" => rgb <= "110110";
					when "11101001110" => rgb <= "110110";
					when "11101001111" => rgb <= "110110";
					when "11101010000" => rgb <= "110110";
					when "11101010001" => rgb <= "110110";
					when "11101010010" => rgb <= "110110";
					when "11101010011" => rgb <= "110110";
					when "11101010100" => rgb <= "110110";
					when "11101010101" => rgb <= "110110";
					when "11101010110" => rgb <= "110110";
					when "11101010111" => rgb <= "110110";
					when "11101011000" => rgb <= "110110";
					when "11101011001" => rgb <= "110110";
					when "11101100000" => rgb <= "110110";
					when "11101100001" => rgb <= "110110";
					when "11101100010" => rgb <= "000000";
					when "11101100011" => rgb <= "000000";
					when "11101100100" => rgb <= "000000";
					when "11101100101" => rgb <= "000000";
					when "11101100110" => rgb <= "000000";
					when "11101100111" => rgb <= "000000";
					when "11101101000" => rgb <= "110110";
					when "11101101001" => rgb <= "110110";
					when "11101101010" => rgb <= "110110";
					when "11101101011" => rgb <= "110110";
					when "11101101100" => rgb <= "110110";
					when "11101101101" => rgb <= "110110";
					when "11101101110" => rgb <= "110110";
					when "11101101111" => rgb <= "110110";
					when "11101110000" => rgb <= "110110";
					when "11101110001" => rgb <= "110110";
					when "11101110010" => rgb <= "110110";
					when "11101110011" => rgb <= "110110";
					when "11101110100" => rgb <= "110110";
					when "11101110101" => rgb <= "110110";
					when "11101110110" => rgb <= "110110";
					when "11101110111" => rgb <= "110110";
					when "11101111000" => rgb <= "110110";
					when "11101111001" => rgb <= "110110";
					when "11110000000" => rgb <= "110110";
					when "11110000001" => rgb <= "110110";
					when "11110000010" => rgb <= "000000";
					when "11110000011" => rgb <= "000000";
					when "11110000100" => rgb <= "000000";
					when "11110000101" => rgb <= "000000";
					when "11110000110" => rgb <= "000000";
					when "11110000111" => rgb <= "000000";
					when "11110001000" => rgb <= "110110";
					when "11110001001" => rgb <= "110110";
					when "11110001010" => rgb <= "110110";
					when "11110001011" => rgb <= "110110";
					when "11110001100" => rgb <= "110110";
					when "11110001101" => rgb <= "110110";
					when "11110001110" => rgb <= "110110";
					when "11110001111" => rgb <= "110110";
					when "11110010000" => rgb <= "110110";
					when "11110010001" => rgb <= "110110";
					when "11110010010" => rgb <= "110110";
					when "11110010011" => rgb <= "110110";
					when "11110010100" => rgb <= "110110";
					when "11110010101" => rgb <= "110110";
					when "11110010110" => rgb <= "110110";
					when "11110010111" => rgb <= "110110";
					when "11110011000" => rgb <= "110110";
					when "11110011001" => rgb <= "110110";
					when "11110100000" => rgb <= "110110";
					when "11110100001" => rgb <= "110110";
					when "11110100010" => rgb <= "000000";
					when "11110100011" => rgb <= "000000";
					when "11110100100" => rgb <= "000000";
					when "11110100101" => rgb <= "000000";
					when "11110100110" => rgb <= "000000";
					when "11110100111" => rgb <= "000000";
					when "11110101000" => rgb <= "110110";
					when "11110101001" => rgb <= "110110";
					when "11110101010" => rgb <= "110110";
					when "11110101011" => rgb <= "110110";
					when "11110101100" => rgb <= "110110";
					when "11110101101" => rgb <= "110110";
					when "11110101110" => rgb <= "110110";
					when "11110101111" => rgb <= "110110";
					when "11110110000" => rgb <= "110110";
					when "11110110001" => rgb <= "110110";
					when "11110110010" => rgb <= "110110";
					when "11110110011" => rgb <= "110110";
					when "11110110100" => rgb <= "110110";
					when "11110110101" => rgb <= "110110";
					when "11110110110" => rgb <= "110110";
					when "11110110111" => rgb <= "110110";
					when "11110111000" => rgb <= "110110";
					when "11110111001" => rgb <= "110110";
					when "11111000000" => rgb <= "110110";
					when "11111000001" => rgb <= "110110";
					when "11111000010" => rgb <= "110110";
					when "11111000011" => rgb <= "110110";
					when "11111000100" => rgb <= "000000";
					when "11111000101" => rgb <= "000000";
					when "11111000110" => rgb <= "000000";
					when "11111000111" => rgb <= "000000";
					when "11111001000" => rgb <= "000000";
					when "11111001001" => rgb <= "000000";
					when "11111001010" => rgb <= "110110";
					when "11111001011" => rgb <= "110110";
					when "11111001100" => rgb <= "110110";
					when "11111001101" => rgb <= "110110";
					when "11111001110" => rgb <= "110110";
					when "11111001111" => rgb <= "110110";
					when "11111010000" => rgb <= "110110";
					when "11111010001" => rgb <= "110110";
					when "11111010010" => rgb <= "110110";
					when "11111010011" => rgb <= "110110";
					when "11111010100" => rgb <= "110110";
					when "11111010101" => rgb <= "110110";
					when "11111010110" => rgb <= "110110";
					when "11111010111" => rgb <= "110110";
					when "11111011000" => rgb <= "110110";
					when "11111011001" => rgb <= "110110";
					when "11111100000" => rgb <= "110110";
					when "11111100001" => rgb <= "110110";
					when "11111100010" => rgb <= "110110";
					when "11111100011" => rgb <= "110110";
					when "11111100100" => rgb <= "000000";
					when "11111100101" => rgb <= "000000";
					when "11111100110" => rgb <= "000000";
					when "11111100111" => rgb <= "000000";
					when "11111101000" => rgb <= "000000";
					when "11111101001" => rgb <= "000000";
					when "11111101010" => rgb <= "110110";
					when "11111101011" => rgb <= "110110";
					when "11111101100" => rgb <= "110110";
					when "11111101101" => rgb <= "110110";
					when "11111101110" => rgb <= "110110";
					when "11111101111" => rgb <= "110110";
					when "11111110000" => rgb <= "110110";
					when "11111110001" => rgb <= "110110";
					when "11111110010" => rgb <= "110110";
					when "11111110011" => rgb <= "110110";
					when "11111110100" => rgb <= "110110";
					when "11111110101" => rgb <= "110110";
					when "11111110110" => rgb <= "110110";
					when "11111110111" => rgb <= "110110";
					when "11111111000" => rgb <= "110110";
					when "11111111001" => rgb <= "110110";
					when others => rgb <= "111111";
		end case;
	end if;
   end process;
   totaladr <= std_logic_vector(yadr) & std_logic_vector(xadr);
end;